//////////////////////////TB_  irq_if ////////////////////////
//DUT interfaces
//////////////////////////////////////////////////////////////////
interface irq_if;

  logic c; 
  logic uc;
  
endinterface: irq_if

