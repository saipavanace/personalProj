
////////////////////////////////////////////////////////////////////////////////
//
// CHI node parameters package
//
////////////////////////////////////////////////////////////////////////////////

package <%=obj.BlockId%>_svt_chi_node_params_pkg;

    `include "<%=obj.BlockId%>_chi_widths.svh"

endpackage : <%=obj.BlockId%>_svt_chi_node_params_pkg
