package dve_seq_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import sv_assert_pkg::*;
  import addr_trans_mgr_pkg::*;
  import dve0_smi_agent_pkg::*;
//  import dve_unit_args_pkg::*;

  `include "dve_coverage_seq.svh"
  `include "dve_cntr.svh"
  `include "dve_seq.svh"
  `include "dve_targt_id_err_seq.svh"
endpackage: dve_seq_pkg
