

parameter integer nACEs       = 1;
parameter integer nACElites   = 0;
parameter integer nAIUs       = 1;
parameter integer nCBIs     = 0;
parameter integer nDCEs       = 1;
parameter integer nDMIs       = 1;
parameter integer vUnitIDAIU0 = 0;
parameter integer vUnitIDAIU1 = 1;
parameter integer vUnitIDAIU2 = 2;
parameter integer vUnitIDAIU3 = 3;
parameter integer vUnitIDDCE  = 4;
parameter integer vUnitIDDMI  = 5;

parameter integer nSFIMasters = nAIUs + nCBIs + nDCEs + nDMIs;
parameter integer nSFISlaves  = nAIUs + nCBIs + nDCEs + nDMIs;

