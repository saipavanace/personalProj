package common_knob_pkg;
    import uvm_pkg::*;
    `include "common_knob_class.svh"
    `include "common_knob_list.svh"
endpackage : common_knob_pkg
