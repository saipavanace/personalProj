// File to control constraints from sequences
//`include "chi_ss_helper_pkg.sv"
// List of all sequence items used in CHI subsys
`include "chi_subsys_base_item.sv"
`include "chi_subsys_snoop_base_item.sv"
`include "chi_subsys_noatomic_item.sv"
`include "chi_subsys_regular_cohexcl_item.sv"
`include "chi_subsys_atomic_compare_item.sv"
`include "chi_subsys_atomic_item.sv"
`include "chi_subsys_regular_item.sv"
`include "chi_subsys_regular_perf_item.sv"
`include "chi_subsys_regular_noncoh_item.sv"
`include "chi_subsys_error_item.sv"
`include "chi_subsys_force_error_item.sv"
`include "chi_subsys_force_snoop_error_item.sv"
`include "chi_subsys_snoop_perf_item.sv"
`include "chi_subsys_regular_error_item.sv"
`include "chi_subsys_snoop_error_item.sv"
`include "chi_subsys_snoop_ptl_resp_item.sv"
`include "chi_subsys_copyback_item.sv"
`include "chi_subsys_nondata_item.sv"
`include "chi_subsys_stash_item.sv"
`include "chi_subsys_connectivity_item.sv"
// List of all sequences used in CHI subsys
`include "chi_subsys_base_seq.sv"
`include "chi_subsys_dvmop_seq.sv"
`include "chi_subsys_mkrdunq_error_seq.sv"
`include "chi_subsys_write_excl_seq.sv"
`include "chi_subsys_comb_wrcmo_seq.sv"
`include "chi_subsys_unsupported_txn_seq.sv"
`include "chi_subsys_atomic_stress_seq.sv"
`include "chi_subsys_stash_stress_seq.sv"
`include "chi_subsys_ip_error_seq.sv"
`include "chi_subsys_random_seq.sv"
`include "chi_subsys_error_seq.sv"
`include "chi_subsys_snp_seq.sv"
`include "chi_subsys_perf_seq.sv"
`include "chi_subsys_random_noncoh_seq.sv"
`include "chi_subsys_random_coherency_seq.sv"
`include "chi_subsys_cmo_seq.sv"
`include "chi_subsys_directed_seq.sv"
`include "chi_subsys_noncoh_seq.sv"
`include "chi_subsys_read_directed_seq.sv"
`include "chi_subsys_directed_noncoh_wr_rd_check_seq.sv"
`include "chi_subsys_multicopy_atomicity_wr_seq.sv"
`include "svt_chi_consumer_seq.svh"
`include "chi_subsys_directed_atomic_self_check_seq.sv"
`include "chi_subsys_directed_coh_wr_rd_check_seq.sv"
`include "chi_subsys_rd_txn_directed_seq.sv"
`include "chi_subsys_coherency_entry_seq.sv"
`include "chi_subsys_directed_snp_resp_seq.sv"
`include "chi_subsys_mkrdunq_seq.sv"
`include "chi_subsys_wrevctorevct_seq.sv"
`include "chi_subsys_directed_atomic_seq.sv"
`include "chi_subsys_owo_writes_seq.sv"
