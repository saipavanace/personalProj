package <%=obj.BlockId%>_trace_debug_env_pkg;
   import uvm_pkg::*;

`include "<%=obj.BlockId%>_trace_debug_env.sv";
endpackage : <%=obj.BlockId%>_trace_debug_env_pkg
