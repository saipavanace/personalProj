
package <%=obj.BlockId%>_axi_slv_mem_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"


import <%=obj.BlockId%>_axi_pkg::*;
import <%=obj.BlockId%>_axi_seq_lib_pkg::*;

`include "<%=obj.BlockId%>_axi_slv_mem_modal.svh"

endpackage: <%=obj.BlockId%>_axi_slv_mem_pkg
