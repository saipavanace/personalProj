package <%=obj.BlockId%>_dirm_pkg;
   import uvm_pkg::*;
`include "uvm_macros.svh"
   import <%=obj.BlockId%>_ConcertoPkg::*;
   
   import addr_trans_mgr_pkg::*;
   
   `include "<%=obj.BlockId%>_dce_dirm_model.svh"     
endpackage 
//
   
   
