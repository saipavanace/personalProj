
class ncore_partial_boot_vseq extends uvm_sequence;
  `uvm_object_utils(ncore_partial_boot_vseq)
  
  
  
  function new(string name = "ncore_partial_boot_vseq");
    super.new(name);
  endfunction: new
  
  virtual task pre_body();
  endtask: pre_body
  
  virtual task body();
    super.body();
      
  
  endtask: body

endclass: ncore_partial_boot_vseq

