////////////////////////////////////////////////////////////////////////////////
//
// Q Channel Agent Package
//
////////////////////////////////////////////////////////////////////////////////
package q_chnl_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "q_chnl_seq_item.svh"
`include "q_chnl_seq.sv"
//`include "q_chnl_if.sv"
`include "q_chnl_agent_config.svh"
`include "q_chnl_driver.svh"
`include "q_chnl_monitor.svh"
`include "q_chnl_sequencer.svh"
`include "q_chnl_agent.svh"

endpackage : q_chnl_agent_pkg
