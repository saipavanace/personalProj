//////////////////////////TB_  IRQ_if ////////////////////////
//DUT interfaces
//////////////////////////////////////////////////////////////////
interface ncore_irq_if;

  wire IRQ_c; 
  wire IRQ_uc;
  
endinterface: ncore_irq_if

