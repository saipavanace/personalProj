

module fsys_config1 (
input 		clk,
input 		reset_n,
input [ 6 : 0]	ioaiuMyId,
output 		awready,
input 		awvalid,
input [ 11 : 0]	awid,
input [ 31 : 0]	awaddr,
input [ 7 : 0]	awlen,
input [ 2 : 0]	awsize,
input [ 1 : 0]	awburst,
input 		awlock,
input [ 3 : 0]	awcache,
input [ 2 : 0]	awprot,
input [ 3 : 0]	awqos,
input [ 11 : 0]	awuser,
input [ 1 : 0]	awdomain,
input [ 2 : 0]	awsnoop,
input [ 1 : 0]	awbar,
output 		wready,
input 		wvalid,
input [ 127 : 0]	wdata,
input [ 15 : 0]	wstrb,
input 		wlast,
input 		bready,
output 		bvalid,
output [ 11 : 0]	bid,
output [ 1 : 0]	bresp,
output 		arready,
input 		arvalid,
input [ 11 : 0]	arid,
input [ 31 : 0]	araddr,
input [ 7 : 0]	arlen,
input [ 2 : 0]	arsize,
input [ 1 : 0]	arburst,
input 		arlock,
input [ 3 : 0]	arcache,
input [ 2 : 0]	arprot,
input [ 3 : 0]	arqos,
input [ 11 : 0]	aruser,
input [ 1 : 0]	ardomain,
input [ 3 : 0]	arsnoop,
input [ 1 : 0]	arbar,
input 		rready,
output 		rvalid,
output [ 11 : 0]	rid,
output [ 127 : 0]	rdata,
output [ 1 : 0]	rresp,
output 		rlast,
output [ 11 : 0]	ruser);



wire  	        io_smi_nd_msg0_tx_ndp_valid;
wire 	        io_smi_nd_msg0_tx_ndp_ready;
wire  [ 7 : 0]	io_smi_nd_msg0_tx_ndp_pbits;
wire  	        io_smi_nd_msg0_tx_ndp_dp_present;
wire  [ 9 : 0]	io_smi_nd_msg0_tx_ndp_target_id;
wire  [ 9 : 0]	io_smi_nd_msg0_tx_ndp_initiator_id;
wire  [ 9 : 0]	io_smi_nd_msg0_tx_ndp_message_id;
wire  [ 7 : 0]	io_smi_nd_msg0_tx_ndp_cm_type;
wire  [ 7 : 0]	io_smi_nd_msg0_tx_ndp_h_prot;
wire  [ 2 : 0]	io_smi_nd_msg0_tx_ndp_t_tier;
wire  [ 2 : 0]	io_smi_nd_msg0_tx_ndp_steering;
wire  [ 2 : 0]	io_smi_nd_msg0_tx_ndp_priority;
wire  [ 2 : 0]	io_smi_nd_msg0_tx_ndp_ql;
wire  [102 : 0]	io_smi_nd_msg0_tx_ndp_body;
wire        	io_smi_nd_msg1_tx_ndp_valid;
wire        	io_smi_nd_msg1_tx_ndp_ready;
wire  [ 7 : 0]	io_smi_nd_msg1_tx_ndp_pbits;
wire  	        io_smi_nd_msg1_tx_ndp_dp_present;
wire  [ 9 : 0]	io_smi_nd_msg1_tx_ndp_target_id;
wire  [ 9 : 0]	io_smi_nd_msg1_tx_ndp_initiator_id;
wire  [ 9 : 0]	io_smi_nd_msg1_tx_ndp_message_id;
wire  [ 7 : 0]	io_smi_nd_msg1_tx_ndp_cm_type;
wire  [ 7 : 0]	io_smi_nd_msg1_tx_ndp_h_prot;
wire  [ 2 : 0]	io_smi_nd_msg1_tx_ndp_t_tier;
wire  [ 2 : 0]	io_smi_nd_msg1_tx_ndp_steering;
wire  [ 2 : 0]	io_smi_nd_msg1_tx_ndp_priority;
wire  [ 2 : 0]	io_smi_nd_msg1_tx_ndp_ql;
wire  [ 102 :0] io_smi_nd_msg1_tx_ndp_body;
wire  	        io_smi_nd_msg2_tx_ndp_valid;
wire 	        io_smi_nd_msg2_tx_ndp_ready;
wire  [ 7 : 0]	io_smi_nd_msg2_tx_ndp_pbits;
wire  	        io_smi_nd_msg2_tx_ndp_dp_present;
wire  [ 2 : 0]	io_smi_nd_msg2_tx_ndp_cdwid;
wire  [ 9 : 0]	io_smi_nd_msg2_tx_ndp_target_id;
wire  [ 9 : 0]	io_smi_nd_msg2_tx_ndp_initiator_id;
wire  [ 9 : 0]	io_smi_nd_msg2_tx_ndp_message_id;
wire  [ 7 : 0]	io_smi_nd_msg2_tx_ndp_cm_type;
wire  [ 7 : 0]	io_smi_nd_msg2_tx_ndp_h_prot;
wire  [ 2 : 0]	io_smi_nd_msg2_tx_ndp_t_tier;
wire  [ 2 : 0]	io_smi_nd_msg2_tx_ndp_steering;
wire  [ 2 : 0]	io_smi_nd_msg2_tx_ndp_priority;
wire  [ 2 : 0]	io_smi_nd_msg2_tx_ndp_ql;
wire  [102 : 0]	io_smi_nd_msg2_tx_ndp_body;
wire        	io_smi_nd_msg2_tx_dp_valid;
wire 	        io_smi_nd_msg2_tx_dp_ready;
wire  	        io_smi_nd_msg2_tx_dp_last;
wire [ 127 : 0] io_smi_nd_msg2_tx_dp_data;
wire  [ 23 : 0] io_smi_nd_msg2_tx_dp_aux;
wire 	        io_smi_nd_msg0_rx_ndp_valid;
wire  	        io_smi_nd_msg0_rx_ndp_ready;
wire [ 7 : 0]	io_smi_nd_msg0_rx_ndp_pbits;
wire 	        io_smi_nd_msg0_rx_ndp_dp_present;
wire [ 9 : 0]	io_smi_nd_msg0_rx_ndp_target_id;
wire [ 9 : 0]	io_smi_nd_msg0_rx_ndp_initiator_id;
wire [ 9 : 0]	io_smi_nd_msg0_rx_ndp_message_id;
wire [ 7 : 0]	io_smi_nd_msg0_rx_ndp_cm_type;
wire [ 7 : 0]	io_smi_nd_msg0_rx_ndp_h_prot;
wire [ 2 : 0]	io_smi_nd_msg0_rx_ndp_t_tier;
wire [ 2 : 0]	io_smi_nd_msg0_rx_ndp_steering;
wire [ 2 : 0]	io_smi_nd_msg0_rx_ndp_priority;
wire [ 2 : 0]	io_smi_nd_msg0_rx_ndp_ql;
wire [ 102 : 0] io_smi_nd_msg0_rx_ndp_body;
wire 	        io_smi_nd_msg1_rx_ndp_valid;
wire         	io_smi_nd_msg1_rx_ndp_ready;
wire [ 7 : 0]	io_smi_nd_msg1_rx_ndp_pbits;
wire 	        io_smi_nd_msg1_rx_ndp_dp_present;
wire [ 9 : 0]	io_smi_nd_msg1_rx_ndp_target_id;
wire [ 9 : 0]	io_smi_nd_msg1_rx_ndp_initiator_id;
wire [ 9 : 0]	io_smi_nd_msg1_rx_ndp_message_id;
wire [ 7 : 0]	io_smi_nd_msg1_rx_ndp_cm_type;
wire [ 7 : 0]	io_smi_nd_msg1_rx_ndp_h_prot;
wire [ 2 : 0]	io_smi_nd_msg1_rx_ndp_t_tier;
wire [ 2 : 0]	io_smi_nd_msg1_rx_ndp_steering;
wire [ 2 : 0]	io_smi_nd_msg1_rx_ndp_priority;
wire [ 2 : 0]	io_smi_nd_msg1_rx_ndp_ql;
wire [102 : 0]	io_smi_nd_msg1_rx_ndp_body;
wire       	    io_smi_nd_msg2_rx_ndp_valid;
wire  	        io_smi_nd_msg2_rx_ndp_ready;
wire [ 7 : 0]	io_smi_nd_msg2_rx_ndp_pbits;
wire 	        io_smi_nd_msg2_rx_ndp_dp_present;
wire [ 2 : 0]	io_smi_nd_msg2_rx_ndp_cdwid;
wire [ 9 : 0]	io_smi_nd_msg2_rx_ndp_target_id;
wire [ 9 : 0]	io_smi_nd_msg2_rx_ndp_initiator_id;
wire [ 9 : 0]	io_smi_nd_msg2_rx_ndp_message_id;
wire [ 7 : 0]	io_smi_nd_msg2_rx_ndp_cm_type;
wire [ 7 : 0]	io_smi_nd_msg2_rx_ndp_h_prot;
wire [ 2 : 0]	io_smi_nd_msg2_rx_ndp_t_tier;
wire [ 2 : 0]	io_smi_nd_msg2_rx_ndp_steering;
wire [ 2 : 0]	io_smi_nd_msg2_rx_ndp_priority;
wire [ 2 : 0]	io_smi_nd_msg2_rx_ndp_ql;
wire [102 : 0]	io_smi_nd_msg2_rx_ndp_body;
wire        	io_smi_nd_msg2_rx_dp_valid;
wire  	        io_smi_nd_msg2_rx_dp_ready;
wire 	        io_smi_nd_msg2_rx_dp_last;
wire [ 127 : 0] io_smi_nd_msg2_rx_dp_data;
wire [ 16 : 0]	io_smi_nd_msg2_rx_dp_aux;

ioaiu_top u_ioaiu(
         .clk(clk),
         .reset_n(reset_n),
         .MyId(ioaiuMyId),
         .awready(awready),
         .awvalid(awvalid),
         .awid(awid),
         .awaddr(awaddr),
         .awlen(awlen),
         .awsize(awsize),
         .awburst(awburst),
         .awlock(awlock),
         .awcache(awcache),
         .awprot(awprot),
         .awqos(awqos),
         .awuser(awuser),
         .awdomain(awdomain),
         .awsnoop(awsnoop),
         .awbar(awbar),
         .wready(wready),
         .wvalid(wvalid),
         .wdata(wdata),
         .wstrb(wstrb),
         .wlast(wlast),
         .bready(bready),
         .bvalid(bvalid),
         .bid(bid),
         .bresp(bresp),
         .arready(arready),
         .arvalid(arvalid),
         .arid(arid),
         .araddr(araddr),
         .arlen(arlen),
         .arsize(arsize),
         .arburst(arburst),
         .arlock(arlock),
         .arcache(arcache),
         .arprot(arprot),
         .arqos(arqos),
         .aruser(aruser),
         .ardomain(ardomain),
         .arsnoop(arsnoop),
         .arbar(arbar),
         .rready(rready),
         .rvalid(rvalid),
         .rid(rid),
         .rdata(rdata),
         .rresp(rresp),
         .rlast(rlast),
         .ruser(ruser),
         .smi_nd_msg0_tx_ndp_valid(io_smi_nd_msg0_tx_ndp_valid),
         .smi_nd_msg0_tx_ndp_ready(io_smi_nd_msg0_tx_ndp_ready),
         .smi_nd_msg0_tx_ndp_pbits(io_smi_nd_msg0_tx_ndp_pbits),
         .smi_nd_msg0_tx_ndp_dp_present(io_smi_nd_msg0_tx_ndp_dp_present),
         .smi_nd_msg0_tx_ndp_target_id(io_smi_nd_msg0_tx_ndp_target_id),
         .smi_nd_msg0_tx_ndp_initiator_id(io_smi_nd_msg0_tx_ndp_initiator_id),
         .smi_nd_msg0_tx_ndp_message_id(io_smi_nd_msg0_tx_ndp_message_id),
         .smi_nd_msg0_tx_ndp_cm_type(io_smi_nd_msg0_tx_ndp_cm_type),
         .smi_nd_msg0_tx_ndp_h_prot(io_smi_nd_msg0_tx_ndp_h_prot),
         .smi_nd_msg0_tx_ndp_t_tier(io_smi_nd_msg0_tx_ndp_t_tier),
         .smi_nd_msg0_tx_ndp_steering(io_smi_nd_msg0_tx_ndp_steering),
         .smi_nd_msg0_tx_ndp_priority(io_smi_nd_msg0_tx_ndp_priority),
         .smi_nd_msg0_tx_ndp_ql(io_smi_nd_msg0_tx_ndp_ql),
         .smi_nd_msg0_tx_ndp_body(io_smi_nd_msg0_tx_ndp_body),
         .smi_nd_msg1_tx_ndp_valid(io_smi_nd_msg1_tx_ndp_valid),
         .smi_nd_msg1_tx_ndp_ready(io_smi_nd_msg1_tx_ndp_ready),
         .smi_nd_msg1_tx_ndp_pbits(io_smi_nd_msg1_tx_ndp_pbits),
         .smi_nd_msg1_tx_ndp_dp_present(io_smi_nd_msg1_tx_ndp_dp_present),
         .smi_nd_msg1_tx_ndp_target_id(io_smi_nd_msg1_tx_ndp_target_id),
         .smi_nd_msg1_tx_ndp_initiator_id(io_smi_nd_msg1_tx_ndp_initiator_id),
         .smi_nd_msg1_tx_ndp_message_id(io_smi_nd_msg1_tx_ndp_message_id),
         .smi_nd_msg1_tx_ndp_cm_type(io_smi_nd_msg1_tx_ndp_cm_type),
         .smi_nd_msg1_tx_ndp_h_prot(io_smi_nd_msg1_tx_ndp_h_prot),
         .smi_nd_msg1_tx_ndp_t_tier(io_smi_nd_msg1_tx_ndp_t_tier),
         .smi_nd_msg1_tx_ndp_steering(io_smi_nd_msg1_tx_ndp_steering),
         .smi_nd_msg1_tx_ndp_priority(io_smi_nd_msg1_tx_ndp_priority),
         .smi_nd_msg1_tx_ndp_ql(io_smi_nd_msg1_tx_ndp_ql),
         .smi_nd_msg1_tx_ndp_body(io_smi_nd_msg1_tx_ndp_body),
         .smi_nd_msg2_tx_ndp_valid(io_smi_nd_msg2_tx_ndp_valid),
         .smi_nd_msg2_tx_ndp_ready(io_smi_nd_msg2_tx_ndp_ready),
         .smi_nd_msg2_tx_ndp_pbits(io_smi_nd_msg2_tx_ndp_pbits),
         .smi_nd_msg2_tx_ndp_dp_present(io_smi_nd_msg2_tx_ndp_dp_present),
         .smi_nd_msg2_tx_ndp_cdwid(io_smi_nd_msg2_tx_ndp_cdwid),
         .smi_nd_msg2_tx_ndp_target_id(io_smi_nd_msg2_tx_ndp_target_id),
         .smi_nd_msg2_tx_ndp_initiator_id(io_smi_nd_msg2_tx_ndp_initiator_id),
         .smi_nd_msg2_tx_ndp_message_id(io_smi_nd_msg2_tx_ndp_message_id),
         .smi_nd_msg2_tx_ndp_cm_type(io_smi_nd_msg2_tx_ndp_cm_type),
         .smi_nd_msg2_tx_ndp_h_prot(io_smi_nd_msg2_tx_ndp_h_prot),
         .smi_nd_msg2_tx_ndp_t_tier(io_smi_nd_msg2_tx_ndp_t_tier),
         .smi_nd_msg2_tx_ndp_steering(io_smi_nd_msg2_tx_ndp_steering),
         .smi_nd_msg2_tx_ndp_priority(io_smi_nd_msg2_tx_ndp_priority),
         .smi_nd_msg2_tx_ndp_ql(io_smi_nd_msg2_tx_ndp_ql),
         .smi_nd_msg2_tx_ndp_body(io_smi_nd_msg2_tx_ndp_body),
         .smi_nd_msg2_tx_dp_valid(io_smi_nd_msg2_tx_dp_valid),
         .smi_nd_msg2_tx_dp_ready(io_smi_nd_msg2_tx_dp_ready),
         .smi_nd_msg2_tx_dp_last(io_smi_nd_msg2_tx_dp_last),
         .smi_nd_msg2_tx_dp_data(io_smi_nd_msg2_tx_dp_data),
         .smi_nd_msg2_tx_dp_aux(io_smi_nd_msg2_tx_dp_aux),
         .smi_nd_msg0_rx_ndp_valid(io_smi_nd_msg0_rx_ndp_valid),
         .smi_nd_msg0_rx_ndp_ready(io_smi_nd_msg0_rx_ndp_ready),
         .smi_nd_msg0_rx_ndp_pbits(io_smi_nd_msg0_rx_ndp_pbits),
         .smi_nd_msg0_rx_ndp_dp_present(io_smi_nd_msg0_rx_ndp_dp_present),
         .smi_nd_msg0_rx_ndp_target_id(io_smi_nd_msg0_rx_ndp_target_id),
         .smi_nd_msg0_rx_ndp_initiator_id(io_smi_nd_msg0_rx_ndp_initiator_id),
         .smi_nd_msg0_rx_ndp_message_id(io_smi_nd_msg0_rx_ndp_message_id),
         .smi_nd_msg0_rx_ndp_cm_type(io_smi_nd_msg0_rx_ndp_cm_type),
         .smi_nd_msg0_rx_ndp_h_prot(io_smi_nd_msg0_rx_ndp_h_prot),
         .smi_nd_msg0_rx_ndp_t_tier(io_smi_nd_msg0_rx_ndp_t_tier),
         .smi_nd_msg0_rx_ndp_steering(io_smi_nd_msg0_rx_ndp_steering),
         .smi_nd_msg0_rx_ndp_priority(io_smi_nd_msg0_rx_ndp_priority),
         .smi_nd_msg0_rx_ndp_ql(io_smi_nd_msg0_rx_ndp_ql),
         .smi_nd_msg0_rx_ndp_body(io_smi_nd_msg0_rx_ndp_body),
         .smi_nd_msg1_rx_ndp_valid(io_smi_nd_msg1_rx_ndp_valid),
         .smi_nd_msg1_rx_ndp_ready(io_smi_nd_msg1_rx_ndp_ready),
         .smi_nd_msg1_rx_ndp_pbits(io_smi_nd_msg1_rx_ndp_pbits),
         .smi_nd_msg1_rx_ndp_dp_present(io_smi_nd_msg1_rx_ndp_dp_present),
         .smi_nd_msg1_rx_ndp_target_id(io_smi_nd_msg1_rx_ndp_target_id),
         .smi_nd_msg1_rx_ndp_initiator_id(io_smi_nd_msg1_rx_ndp_initiator_id),
         .smi_nd_msg1_rx_ndp_message_id(io_smi_nd_msg1_rx_ndp_message_id),
         .smi_nd_msg1_rx_ndp_cm_type(io_smi_nd_msg1_rx_ndp_cm_type),
         .smi_nd_msg1_rx_ndp_h_prot(io_smi_nd_msg1_rx_ndp_h_prot),
         .smi_nd_msg1_rx_ndp_t_tier(io_smi_nd_msg1_rx_ndp_t_tier),
         .smi_nd_msg1_rx_ndp_steering(io_smi_nd_msg1_rx_ndp_steering),
         .smi_nd_msg1_rx_ndp_priority(io_smi_nd_msg1_rx_ndp_priority),
         .smi_nd_msg1_rx_ndp_ql(io_smi_nd_msg1_rx_ndp_ql),
         .smi_nd_msg1_rx_ndp_body(io_smi_nd_msg1_rx_ndp_body),
         .smi_nd_msg2_rx_ndp_valid(io_smi_nd_msg2_rx_ndp_valid),
         .smi_nd_msg2_rx_ndp_ready(io_smi_nd_msg2_rx_ndp_ready),
         .smi_nd_msg2_rx_ndp_pbits(io_smi_nd_msg2_rx_ndp_pbits),
         .smi_nd_msg2_rx_ndp_dp_present(io_smi_nd_msg2_rx_ndp_dp_present),
         .smi_nd_msg2_rx_ndp_cdwid(io_smi_nd_msg2_rx_ndp_cdwid),
         .smi_nd_msg2_rx_ndp_target_id(io_smi_nd_msg2_rx_ndp_target_id),
         .smi_nd_msg2_rx_ndp_message_id(io_smi_nd_msg2_rx_ndp_message_id),
         .smi_nd_msg2_rx_ndp_cm_type(io_smi_nd_msg2_rx_ndp_cm_type),
         .smi_nd_msg2_rx_ndp_h_prot(io_smi_nd_msg2_rx_ndp_h_prot),
         .smi_nd_msg2_rx_ndp_t_tier(io_smi_nd_msg2_rx_ndp_t_tier),
         .smi_nd_msg2_rx_ndp_steering(io_smi_nd_msg2_rx_ndp_steering),
         .smi_nd_msg2_rx_ndp_priority(io_smi_nd_msg2_rx_ndp_priority),
         .smi_nd_msg2_rx_ndp_ql(io_smi_nd_msg2_rx_ndp_ql),
         .smi_nd_msg2_rx_ndp_body(io_smi_nd_msg2_rx_ndp_body),
         .smi_nd_msg2_rx_dp_valid(io_smi_nd_msg2_rx_dp_valid),
         .smi_nd_msg2_rx_dp_ready(io_smi_nd_msg2_rx_dp_ready),
         .smi_nd_msg2_rx_dp_last(io_smi_nd_msg2_rx_dp_last),
         .smi_nd_msg2_rx_dp_data(io_smi_nd_msg2_rx_dp_data),
         .smi_nd_msg2_rx_dp_aux(io_smi_nd_msg2_rx_dp_aux),
         .smi_nd_msg2_rx_ndp_initiator_id(io_smi_nd_msg2_rx_ndp_initiator_id)
);

top_wrapper lagato (
 .a_clk(clk),
 .a_reset_n(reset_n),
 .ismi0_valid(io_smi_nd_msg0_tx_ndp_valid),
 .ismi0_ready(io_smi_nd_msg0_tx_ndp_ready),
 .ismi0_targ_id(io_smi_nd_msg0_tx_ndp_target_id),
 .ismi0_route('b0),
 .ismi0_src_id(io_smi_nd_msg0_tx_ndp_initiator_id),
 .ismi0_tier(io_smi_nd_msg0_tx_ndp_t_tier),
 .ismi0_dp_present(io_smi_nd_msg0_tx_ndp_dp_present),
 .ismi0_ndp_len(io_smi_nd_msg0_tx_ndp_pbits),
 .ismi0_ndp(io_smi_nd_msg0_tx_ndp_body),
 .ismi0_msg_type(io_smi_nd_msg0_tx_ndp_cm_type),
 .ismi0_msg_id(io_smi_nd_msg0_tx_ndp_message_id),
 .ismi0_deassert_ready('b0),
 .ismi0_dp_valid('b0),
// .ismi0_dp_ready,
// .ismi0_dp_last,
// .ismi0_dp_data,
// .ismi0_dp_user,
 .ismi1_valid(io_smi_nd_msg1_tx_ndp_valid),
 .ismi1_ready(io_smi_nd_msg1_tx_ndp_ready),
 .ismi1_targ_id(io_smi_nd_msg1_tx_ndp_target_id),
 .ismi1_route('b0),
 .ismi1_src_id(io_smi_nd_msg1_tx_ndp_initiator_id),
 .ismi1_tier(io_smi_nd_msg1_tx_ndp_t_tier),
 .ismi1_dp_present(io_smi_nd_msg1_tx_ndp_dp_present),
 .ismi1_ndp_len(io_smi_nd_msg1_tx_ndp_pbits),
 .ismi1_ndp(io_smi_nd_msg1_tx_ndp_body),
 .ismi1_msg_type(io_smi_nd_msg1_tx_ndp_cm_type),
 .ismi1_msg_id(io_smi_nd_msg1_tx_ndp_message_id),
 .ismi1_deassert_ready('b0),
 .ismi1_dp_valid('b0),
// .ismi1_dp_ready,
// .ismi1_dp_last,
// .ismi1_dp_data,
// .ismi1_dp_user,
 .ismi2_valid(io_smi_nd_msg2_tx_ndp_valid),
 .ismi2_ready(io_smi_nd_msg2_tx_ndp_ready),
 .ismi2_targ_id(io_smi_nd_msg2_tx_ndp_target_id),
 .ismi2_route('b0),
 .ismi2_src_id(io_smi_nd_msg2_tx_ndp_initiator_id),
 .ismi2_tier(io_smi_nd_msg2_tx_ndp_t_tier),
 .ismi2_dp_present(io_smi_nd_msg2_tx_ndp_dp_present),
 .ismi2_ndp_len(io_smi_nd_msg2_tx_ndp_h_prot),
 .ismi2_ndp(io_smi_nd_msg2_tx_ndp_body),
 .ismi2_msg_type(io_smi_nd_msg2_tx_ndp_cm_type),
 .ismi2_msg_id(io_smi_nd_msg2_tx_ndp_message_id),
 .ismi2_deassert_ready('b0),
 .ismi2_dp_valid(io_smi_nd_msg2_tx_dp_valid),
 .ismi2_dp_ready(io_smi_nd_msg2_tx_dp_ready),
 .ismi2_dp_last(io_smi_nd_msg2_tx_dp_last),
 .ismi2_dp_data(io_smi_nd_msg2_tx_dp_data),
 .ismi2_dp_user(io_smi_nd_msg2_tx_dp_aux),
 .ismi3_valid('b0),
// .ismi3_ready,
// .ismi3_targ_id,
// .ismi3_route,
// .ismi3_src_id,
// .ismi3_tier,
// .ismi3_dp_present,
// .ismi3_ndp_len,
// .ismi3_ndp,
// .ismi3_msg_type,
// .ismi3_msg_id,
// .ismi3_deassert_ready,
 .ismi3_dp_valid('b0),
// .ismi3_dp_ready,
// .ismi3_dp_last,
// .ismi3_dp_data,
// .ismi3_dp_user,
 .ismi4_valid('b0),
// .ismi4_ready,
// .ismi4_targ_id,
// .ismi4_route,
// .ismi4_src_id,
// .ismi4_tier,
// .ismi4_dp_present,
// .ismi4_ndp_len,
// .ismi4_ndp,
// .ismi4_msg_type,
// .ismi4_msg_id,
// .ismi4_deassert_ready,
 .ismi4_dp_valid('b0),
// .ismi4_dp_ready,
// .ismi4_dp_last,
// .ismi4_dp_data,
// .ismi4_dp_user,
 .ismi5_valid('b0),
// .ismi5_ready,
// .ismi5_targ_id,
// .ismi5_route,
// .ismi5_src_id,
// .ismi5_tier,
// .ismi5_dp_present,
// .ismi5_ndp_len,
// .ismi5_ndp,
// .ismi5_msg_type,
// .ismi5_msg_id,
// .ismi5_deassert_ready,
 .ismi5_dp_valid('b0),
// .ismi5_dp_ready,
// .ismi5_dp_last,
// .ismi5_dp_data,
// .ismi5_dp_user,
 .ismi6_valid('b0),
// .ismi6_ready,
// .ismi6_targ_id,
// .ismi6_route,
// .ismi6_src_id,
// .ismi6_tier,
// .ismi6_dp_present,
// .ismi6_ndp_len,
// .ismi6_ndp,
// .ismi6_msg_type,
// .ismi6_msg_id,
// .ismi6_deassert_ready,
 .ismi6_dp_valid('b0),
// .ismi6_dp_ready,
// .ismi6_dp_last,
// .ismi6_dp_data,
// .ismi6_dp_user,
 .ismi7_valid('b0),
// .ismi7_ready,
// .ismi7_targ_id,
// .ismi7_route,
// .ismi7_src_id,
// .ismi7_tier,
// .ismi7_dp_present,
// .ismi7_ndp_len,
// .ismi7_ndp,
// .ismi7_msg_type,
// .ismi7_msg_id,
// .ismi7_deassert_ready,
 .ismi7_dp_valid('b0),
// .ismi7_dp_ready,
// .ismi7_dp_last,
// .ismi7_dp_data,
// .ismi7_dp_user,
 .ismi8_valid('b0),
// .ismi8_ready,
// .ismi8_targ_id,
// .ismi8_route,
// .ismi8_src_id,
// .ismi8_tier,
// .ismi8_dp_present,
// .ismi8_ndp_len,
// .ismi8_ndp,
// .ismi8_msg_type,
// .ismi8_msg_id,
// .ismi8_deassert_ready,
 .ismi8_dp_valid('b0),
// .ismi8_dp_ready,
// .ismi8_dp_last,
// .ismi8_dp_data,
// .ismi8_dp_user,
 .ismi9_valid('b0),
// .ismi9_ready,
// .ismi9_targ_id,
// .ismi9_route,
// .ismi9_src_id,
// .ismi9_tier,
// .ismi9_dp_present,
// .ismi9_ndp_len,
// .ismi9_ndp,
// .ismi9_msg_type,
// .ismi9_msg_id,
// .ismi9_deassert_ready,
 .ismi9_dp_valid('b0),
// .ismi9_dp_ready,
// .ismi9_dp_last,
// .ismi9_dp_data,
// .ismi9_dp_user,
 .ismi10_valid('b0),
// .ismi10_ready,
// .ismi10_targ_id,
// .ismi10_route,
// .ismi10_src_id,
// .ismi10_tier,
// .ismi10_dp_present,
// .ismi10_ndp_len,
// .ismi10_ndp,
// .ismi10_msg_type,
// .ismi10_msg_id,
// .ismi10_deassert_ready,
 .ismi10_dp_valid('b0),
// .ismi10_dp_ready,
// .ismi10_dp_last,
// .ismi10_dp_data,
// .ismi10_dp_user,
 .ismi11_valid('b0),
// .ismi11_ready,
// .ismi11_targ_id,
// .ismi11_route,
// .ismi11_src_id,
// .ismi11_tier,
// .ismi11_dp_present,
// .ismi11_ndp_len,
// .ismi11_ndp,
// .ismi11_msg_type,
// .ismi11_msg_id,
// .ismi11_deassert_ready,
 .ismi11_dp_valid('b0),
// .ismi11_dp_ready,
// .ismi11_dp_last,
// .ismi11_dp_data,
// .ismi11_dp_user,
 .ismi12_valid('b0),
// .ismi12_ready,
// .ismi12_targ_id,
// .ismi12_route,
// .ismi12_src_id,
// .ismi12_tier,
// .ismi12_dp_present,
// .ismi12_ndp_len,
// .ismi12_ndp,
// .ismi12_msg_type,
// .ismi12_msg_id,
// .ismi12_deassert_ready,
 .ismi12_dp_valid('b0),
// .ismi12_dp_ready,
// .ismi12_dp_last,
// .ismi12_dp_data,
// .ismi12_dp_user,
 .ismi13_valid('b0),
// .ismi13_ready,
// .ismi13_targ_id,
// .ismi13_route,
// .ismi13_src_id,
// .ismi13_tier,
// .ismi13_dp_present,
// .ismi13_ndp_len,
// .ismi13_ndp,
// .ismi13_msg_type,
// .ismi13_msg_id,
// .ismi13_deassert_ready,
 .ismi13_dp_valid('b0),
// .ismi13_dp_ready,
// .ismi13_dp_last,
// .ismi13_dp_data,
// .ismi13_dp_user,
 .ismi14_valid('b0),
// .ismi14_ready,
// .ismi14_targ_id,
// .ismi14_route,
// .ismi14_src_id,
// .ismi14_tier,
// .ismi14_dp_present,
// .ismi14_ndp_len,
// .ismi14_ndp,
// .ismi14_msg_type,
// .ismi14_msg_id,
// .ismi14_deassert_ready,
 .ismi14_dp_valid('b0),
// .ismi14_dp_ready,
// .ismi14_dp_last,
// .ismi14_dp_data,
// .ismi14_dp_user,
 .ismi15_valid('b0),
// .ismi15_ready,
// .ismi15_targ_id,
// .ismi15_route,
// .ismi15_src_id,
// .ismi15_tier,
// .ismi15_dp_present,
// .ismi15_ndp_len,
// .ismi15_ndp,
// .ismi15_msg_type,
// .ismi15_msg_id,
// .ismi15_deassert_ready,
 .ismi15_dp_valid('b0),
// .ismi15_dp_ready,
// .ismi15_dp_last,
// .ismi15_dp_data,
// .ismi15_dp_user,
 .osmi0_valid(io_smi_nd_msg0_rx_ndp_valid),
 .osmi0_ready(io_smi_nd_msg0_rx_ndp_ready),
 .osmi0_targ_id(io_smi_nd_msg0_rx_ndp_target_id),
 .osmi0_src_id(io_smi_nd_msg0_rx_ndp_initiator_id),
 .osmi0_tier(io_smi_nd_msg0_rx_ndp_t_tier),
 .osmi0_dp_present(io_smi_nd_msg0_rx_ndp_dp_present),
 .osmi0_ndp_len(io_smi_nd_msg0_rx_ndp_pbits),
 .osmi0_ndp(io_smi_nd_msg0_rx_ndp_body),
 .osmi0_msg_type(io_smi_nd_msg0_rx_ndp_cm_type),
 .osmi0_msg_id(io_smi_nd_msg0_rx_ndp_message_id),
// .osmi0_dp_valid,
 .osmi0_dp_ready('b0),
// .osmi0_dp_last,
// .osmi0_dp_data,
// .osmi0_dp_user,
 .osmi1_valid(io_smi_nd_msg1_rx_ndp_valid),
 .osmi1_ready(io_smi_nd_msg1_rx_ndp_ready),
 .osmi1_targ_id(io_smi_nd_msg1_rx_ndp_target_id),
 .osmi1_src_id(io_smi_nd_msg1_rx_ndp_initiator_id),
 .osmi1_tier(io_smi_nd_msg1_rx_ndp_t_tier),
 .osmi1_dp_present(io_smi_nd_msg1_rx_ndp_dp_present),
 .osmi1_ndp_len(io_smi_nd_msg1_rx_ndp_pbits),
 .osmi1_ndp(io_smi_nd_msg1_rx_ndp_body),
 .osmi1_msg_type(io_smi_nd_msg1_rx_ndp_cm_type),
 .osmi1_msg_id(io_smi_nd_msg1_rx_ndp_message_id),
// .osmi1_dp_valid,
 .osmi1_dp_ready('b0),
// .osmi1_dp_last,
// .osmi1_dp_data,
// .osmi1_dp_user,
 .osmi2_valid(io_smi_nd_msg2_rx_ndp_valid),
 .osmi2_ready(io_smi_nd_msg2_rx_ndp_ready),
 .osmi2_targ_id(io_smi_nd_msg2_rx_ndp_target_id),
 .osmi2_src_id(io_smi_nd_msg2_rx_ndp_initiator_id),
 .osmi2_tier(io_smi_nd_msg2_rx_ndp_t_tier),
 .osmi2_dp_present(io_smi_nd_msg2_rx_ndp_dp_present),
 .osmi2_ndp_len(io_smi_nd_msg2_rx_ndp_pbits),
 .osmi2_ndp(io_smi_nd_msg2_rx_ndp_body),
 .osmi2_msg_type(io_smi_nd_msg2_rx_ndp_cm_type),
 .osmi2_msg_id(io_smi_nd_msg2_rx_ndp_message_id),
 .osmi2_dp_valid(io_smi_nd_msg2_rx_dp_valid),
 .osmi2_dp_ready(io_smi_nd_msg2_rx_dp_ready),
 .osmi2_dp_last(io_smi_nd_msg2_rx_dp_last),
 .osmi2_dp_data(io_smi_nd_msg2_rx_dp_data),
 .osmi2_dp_user(io_smi_nd_msg2_rx_dp_aux),
// .osmi3_valid,
 .osmi3_ready('b1),
// .osmi3_targ_id,
// .osmi3_src_id,
// .osmi3_tier,
// .osmi3_dp_present,
// .osmi3_ndp_len,
// .osmi3_ndp,
// .osmi3_msg_type,
// .osmi3_msg_id,
// .osmi3_dp_valid,
 .osmi3_dp_ready('b1),
// .osmi3_dp_last,
// .osmi3_dp_data,
// .osmi3_dp_user,
// .osmi4_valid,
 .osmi4_ready('b1),
// .osmi4_targ_id,
// .osmi4_src_id,
// .osmi4_tier,
// .osmi4_dp_present,
// .osmi4_ndp_len,
// .osmi4_ndp,
// .osmi4_msg_type,
// .osmi4_msg_id,
// .osmi4_dp_valid,
 .osmi4_dp_ready('b1),
// .osmi4_dp_last,
// .osmi4_dp_data,
// .osmi4_dp_user,
// .osmi5_valid,
 .osmi5_ready('b1),
// .osmi5_targ_id,
// .osmi5_src_id,
// .osmi5_tier,
// .osmi5_dp_present,
// .osmi5_ndp_len,
// .osmi5_ndp,
// .osmi5_msg_type,
// .osmi5_msg_id,
// .osmi5_dp_valid,
 .osmi5_dp_ready('b1),
// .osmi5_dp_last,
// .osmi5_dp_data,
// .osmi5_dp_user,
// .osmi6_valid,
 .osmi6_ready('b1),
// .osmi6_targ_id,
// .osmi6_src_id,
// .osmi6_tier,
// .osmi6_dp_present,
// .osmi6_ndp_len,
// .osmi6_ndp,
// .osmi6_msg_type,
// .osmi6_msg_id,
// .osmi6_dp_valid,
 .osmi6_dp_ready('b1),
// .osmi6_dp_last,
// .osmi6_dp_data,
// .osmi6_dp_user,
// .osmi7_valid,
 .osmi7_ready('b1),
// .osmi7_targ_id,
// .osmi7_src_id,
// .osmi7_tier,
// .osmi7_dp_present,
// .osmi7_ndp_len,
// .osmi7_ndp,
// .osmi7_msg_type,
// .osmi7_msg_id,
// .osmi7_dp_valid,
 .osmi7_dp_ready('b1),
// .osmi7_dp_last,
// .osmi7_dp_data,
// .osmi7_dp_user,
// .osmi8_valid,
 .osmi8_ready('b1),
// .osmi8_targ_id,
// .osmi8_src_id,
// .osmi8_tier,
// .osmi8_dp_present,
// .osmi8_ndp_len,
// .osmi8_ndp,
// .osmi8_msg_type,
// .osmi8_msg_id,
// .osmi8_dp_valid,
 .osmi8_dp_ready('b1),
// .osmi8_dp_last,
// .osmi8_dp_data,
// .osmi8_dp_user,
// .osmi9_valid,
 .osmi9_ready('b1),
// .osmi9_targ_id,
// .osmi9_src_id,
// .osmi9_tier,
// .osmi9_dp_present,
// .osmi9_ndp_len,
// .osmi9_ndp,
// .osmi9_msg_type,
// .osmi9_msg_id,
// .osmi9_dp_valid,
 .osmi9_dp_ready('b1),
// .osmi9_dp_last,
// .osmi9_dp_data,
// .osmi9_dp_user,
// .osmi10_valid,
 .osmi10_ready('b1),
// .osmi10_targ_id,
// .osmi10_src_id,
// .osmi10_tier,
// .osmi10_dp_present,
// .osmi10_ndp_len,
// .osmi10_ndp,
// .osmi10_msg_type,
// .osmi10_msg_id,
// .osmi10_dp_valid,
 .osmi10_dp_ready('b1),
// .osmi10_dp_last,
// .osmi10_dp_data,
// .osmi10_dp_user,
// .osmi11_valid,
 .osmi11_ready('b1),
// .osmi11_targ_id,
// .osmi11_src_id,
// .osmi11_tier,
// .osmi11_dp_present,
// .osmi11_ndp_len,
// .osmi11_ndp,
// .osmi11_msg_type,
// .osmi11_msg_id,
// .osmi11_dp_valid,
 .osmi11_dp_ready('b1),
// .osmi11_dp_last,
// .osmi11_dp_data,
// .osmi11_dp_user,
// .osmi12_valid,
 .osmi12_ready('b1),
// .osmi12_targ_id,
// .osmi12_src_id,
// .osmi12_tier,
// .osmi12_dp_present,
// .osmi12_ndp_len,
// .osmi12_ndp,
// .osmi12_msg_type,
// .osmi12_msg_id,
// .osmi12_dp_valid,
 .osmi12_dp_ready('b1),
// .osmi12_dp_last,
// .osmi12_dp_data,
// .osmi12_dp_user,
// .osmi13_valid,
 .osmi13_ready('b1),
// .osmi13_targ_id,
// .osmi13_src_id,
// .osmi13_tier,
// .osmi13_dp_present,
// .osmi13_ndp_len,
// .osmi13_ndp,
// .osmi13_msg_type,
// .osmi13_msg_id,
// .osmi13_dp_valid,
 .osmi13_dp_ready('b1),
// .osmi13_dp_last,
// .osmi13_dp_data,
// .osmi13_dp_user,
// .osmi14_valid,
 .osmi14_ready('b1),
// .osmi14_targ_id,
// .osmi14_src_id,
// .osmi14_tier,
// .osmi14_dp_present,
// .osmi14_ndp_len,
// .osmi14_ndp,
// .osmi14_msg_type,
// .osmi14_msg_id,
// .osmi14_dp_valid,
 .osmi14_dp_ready('b1),
// .osmi14_dp_last,
// .osmi14_dp_data,
// .osmi14_dp_user,
// .osmi15_valid,
 .osmi15_ready('b1),
// .osmi15_targ_id,
// .osmi15_src_id,
// .osmi15_tier,
// .osmi15_dp_present,
// .osmi15_ndp_len,
// .osmi15_ndp,
// .osmi15_msg_type,
// .osmi15_msg_id,
// .osmi15_dp_valid,
 .osmi15_dp_ready('b1)
// .osmi15_dp_last,
// .osmi15_dp_data,
// .osmi15_dp_user 
);

endmodule
