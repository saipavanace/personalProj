`ifndef GUARD_IOAIU_AXI_ACE_MASTER_BASE_VIRTUAL_SEQUENCE_SVH
`define GUARD_IOAIU_AXI_ACE_MASTER_BASE_VIRTUAL_SEQUENCE_SVH

/** Base class from which all ACE basic level sequences will be extended. */
class ioaiu_axi_ace_master_base_virtual_sequence extends svt_axi_ace_master_base_virtual_sequence;
  
  svt_axi_ace_master_base_sequence  coherent_seq;

  ioaiu_axi_ace_master_base_virtual_sequence_controls vseq_controls;
 
  /** Represents the master port from which the sequence will be initiated. */ 
  rand int unsigned port_id; 

  /** Represents the length of the sequence. */
  rand int unsigned sequence_length = 10;

  /** Indicates if this sequence is valid on an ACE port */
  protected bit is_seq_valid_on_ace_port = 1;

  /** Indicates if this sequence is valid on an ACE-Lite port */
  protected bit is_seq_valid_on_ace_lite_port = 1;

  /**
    * The start address for the address range for transactions generated by this
    * sequence. Applicable only for extended sequences where it is specified
    * that start_addr can be provided through uvm_config_db. Typically 
    * applicable only for sequential access sequences.
    */
  bit[`SVT_AXI_ADDR_WIDTH-1:0] start_addr = 0;


  /** Indicates if start_addr has been passed through uvm_config_db, or is directly set */
  bit status_start_addr = 0;
  
  /** If this bit is set to one, transactions are sent to sequential addresses
    * If low, transactions are sent to random addresses
    */
  bit addr_mode_select =0;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer) 

  `svt_xvm_object_utils(ioaiu_axi_ace_master_base_virtual_sequence)

    /** Constrain the sequence length to a reasonable value */
  constraint reasonable_sequence_length {
    sequence_length <= 1000;
  }
   

  function new(string name = "ioaiu_axi_ace_master_base_virtual_sequence");
    super.new(name);
  endfunction

  virtual task pre_body();
    bit status;
    super.pre_body();
    raise_phase_objection();

    status = uvm_config_db#(ioaiu_axi_ace_master_base_virtual_sequence_controls)::get(null, get_full_name(), "vseq_controls", vseq_controls);
    if(status == 0) begin
        `uvm_error("body",$sformatf("vseq_controls of Type=ioaiu_axi_ace_master_base_virtual_sequence_controls is not set properly through uvm_config_db"))
    end
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "sequence_length", sequence_length);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "port_id", port_id);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "addr_mode_select",addr_mode_select );
 
    // If start_addr is already set directly, do not override the status based on whether it was passed
    // through uvm_config_db or not.
    if (!status_start_addr)
      status_start_addr = uvm_config_db#(bit[`SVT_AXI_ADDR_WIDTH-1:0])::get(null, get_full_name(), "start_addr",start_addr);
    
    `svt_xvm_debug("body", $sformatf("port_id is 'd%0d as a result of %0s.", port_id, status ? "config DB" : "randomization"));
    `svt_xvm_debug("body", $sformatf("start_addr is 'h%0h as a result of %0s.", start_addr, status_start_addr ? "config DB" : "randomization"));
  endtask

 /** Drop objection */
  virtual task post_body();
    drop_phase_objection();
  endtask: post_body

  task send_coherent_transactions(svt_axi_transaction::coherent_xact_type_enum master_xact_type ,bit init_cachelines);
    `svt_xvm_create_on(coherent_seq, p_sequencer.master_sequencer[port_id])    
    coherent_seq.assign_xact_weights(master_xact_type);
    coherent_seq.initialize_cachelines = init_cachelines ;
    void'(coherent_seq.randomize with {use_directed_addr == 0;sequence_length==local::sequence_length;});
    coherent_seq.start(p_sequencer.master_sequencer[port_id]); 
  endtask

`ifdef SVT_ACE5_ENABLE
  task send_cmo_on_write_transactions(svt_axi_transaction::coherent_xact_type_enum master_xact_type , svt_axi_transaction::cmo_on_write_xact_type_enum master_cmo_xact_type,bit init_cachelines,bit use_directed_domain_type, svt_axi_transaction::xact_shareability_domain_enum directed_domain_type);
    `svt_xvm_create_on(coherent_seq, p_sequencer.master_sequencer[port_id])    
    coherent_seq.assign_xact_weights(master_xact_type);
    coherent_seq.assign_cmo_on_write_xact_weights(master_cmo_xact_type);
    if(!addr_mode_select)
       coherent_seq.addr_mode = svt_axi_ace_master_base_sequence::RANDOM_ADDR_MODE;
    else 
       coherent_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
    if (use_directed_domain_type) begin
      coherent_seq.use_directed_domain_type = 1;
      coherent_seq.directed_domain_type = directed_domain_type;
    end
    
    if (status_start_addr) begin
      coherent_seq.status_start_addr = 1;
      coherent_seq.start_addr = start_addr;
    end
    
    coherent_seq.initialize_cachelines = init_cachelines ;
    void'(coherent_seq.randomize with {use_directed_addr == 0;sequence_length==local::sequence_length;});
    coherent_seq.start(p_sequencer.master_sequencer[port_id]); 
  endtask
`endif

  virtual function bit is_supported(svt_configuration cfg , bit silent = 0);
    bit is_port_ace = 0;
    bit is_port_ace_lite = 0;
    `svt_xvm_debug("is_supported",$sformatf("calling is_supported")); 
    if (port_id inside {ace_ports})
      is_port_ace = 1;
    else if (port_id inside {ace_lite_ports})
      is_port_ace_lite = 1;

    if (is_seq_valid_on_ace_port) begin
      if (ace_ports.size()) 
        if (is_port_ace)
          is_supported = 1;
    end
    if (is_seq_valid_on_ace_lite_port) begin
      if (ace_lite_ports.size()) 
        if (is_port_ace_lite)
          is_supported = 1;
    end
    if (!is_supported) begin
      if (is_seq_valid_on_ace_port && is_seq_valid_on_ace_lite_port) begin
        `svt_xvm_note("is_supported", $sformatf("port_id('d%0d) is not valid for this sequence. Please ensure  the following: \n\
                                                 svt_axi_port_configuration::axi_interface_type = svt_axi_port_configuration::AXI_ACE or svt_axi_port_configuration::ACE_LITE\n\
                                                 svt_axi_port_configuration::is_active = 1 \n\
                                                 svt_axi_system_configuration::participating_masters[<master>] = 1", port_id));
      end
      else if (is_seq_valid_on_ace_port) begin
        `svt_xvm_note("is_supported", $sformatf("port_id('d%0d) is not valid for this sequence. Please ensure  the following: \n\
                                                 svt_axi_port_configuration::axi_interface_type = svt_axi_port_configuration::AXI_ACE\n\
                                                 svt_axi_port_configuration::is_active = 1 \n\
                                                 svt_axi_system_configuration::participating_masters[<master>] = 1", port_id));
      end
      else if (is_seq_valid_on_ace_lite_port) begin
        `svt_xvm_note("is_supported", $sformatf("port_id('d%0d) is not valid for this sequence. Please ensure  the following: \n\
                                                 svt_axi_port_configuration::axi_interface_type = svt_axi_port_configuration::ACE_LITE\n\
                                                 svt_axi_port_configuration::is_active = 1 \n\
                                                 svt_axi_system_configuration::participating_masters[<master>] = 1", port_id));
      end
    end
    `svt_xvm_debug("is_supported",$sformatf("is_supported = 'd%0d",is_supported)); 
  endfunction

endclass    
 

`endif // `ifndef GUARD_IOAIU_AXI_ACE_MASTER_BASE_VIRTUAL_SEQUENCE_SVH
