// Library of all virtual sequences used in IO Subsystem
`include "io_subsys_snps_base_vseq.svh"
`include "io_subsys_snps_vseq.svh"
`include "io_subsys_snps_pcie_vseq.svh"
`include "io_subsys_stash_stress_vseq.svh"
`include "io_subsys_directed_noncoh_wr_rd_check_vseq.svh"
`include "io_subsys_directed_atomic_self_check_vseq.svh"
`include "io_subsys_directed_coh_wr_rd_check_vseq.svh"
`include "io_subsys_directed_rd_ncaiu_to_all_dmis_noncoh_stress_vseq.svh"
`include "io_subsys_inhouse_base_vseq.svh"
`include "io_subsys_inhouse_vseq.svh"
`include "io_subsys_vseq.svh"
