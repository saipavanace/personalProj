`ifdef USE_VIP_SNPS
   import uvm_pkg::*;
   `include "uvm_macros.svh"
   import svt_uvm_pkg::*;
   import svt_axi_uvm_pkg::*;
`endif
