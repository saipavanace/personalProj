
package <%=obj.BlockId%>_resetPkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "<%=obj.BlockId%>_reset_monitor.svh"

endpackage: <%=obj.BlockId%>_resetPkg
