
package <%=obj.BlockId%>_reset_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

import <%=obj.BlockId%>_ConcertoPkg::*;

`include "<%=obj.BlockId%>_reset_monitor.svh"

endpackage: <%=obj.BlockId%>_reset_pkg
