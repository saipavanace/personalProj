`ifndef DMI_CONFIG_INFO_SV
`define DMI_CONFIG_INFO_SV
`endif
