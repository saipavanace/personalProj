//
// SFI Parameters
//
<% if (obj.testBench == "emu" ) { %>

typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPPOISION-1:0]      <%=obj.BlockId%>_probe_ccp_data_poision_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPDATA-1:0]         <%=obj.BlockId%>_probe_ccp_ctrlwr_data_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_ctrlwr_vld_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPBYTEEN-1:0]       <%=obj.BlockId%>_probe_ccp_ctrlwr_byten_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPBEAT-1:0]         <%=obj.BlockId%>_probe_ccp_ctrlwr_beatn_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_ctrlwr_last_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cachewr_rdy_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_ctrlfilldata_vld_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPDATA-1:0]         <%=obj.BlockId%>_probe_ccp_ctrlfill_data_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPFILLID-1:0]       <%=obj.BlockId%>_probe_ccp_ctrlfilldata_Id_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPADDR-1:0]         <%=obj.BlockId%>_probe_ccp_ctrlfilldata_addr_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPWAYS-1:0]         <%=obj.BlockId%>_probe_ccp_ctrlfilldata_wayn_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPBEAT-1:0]         <%=obj.BlockId%>_probe_ccp_ctrlfilldata_beatn_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPBYTEEN-1:0]       <%=obj.BlockId%>_probe_ccp_ctrlfilldata_byten_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_ctrlfilldata_last_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cachefilldata_rdy_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_ctrlfill_vld_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPADDR-1:0]         <%=obj.BlockId%>_probe_ccp_ctrlfill_addr_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPWAYS-1:0]         <%=obj.BlockId%>_probe_ccp_ctrlfill_wayn_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPSECURITY-1:0]     <%=obj.BlockId%>_probe_ccp_ctrlfill_security_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPCACHESTATE-1:0]   <%=obj.BlockId%>_probe_ccp_ctrlfill_state_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cachefill_rdy_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPFILLDONEID-1:0]   <%=obj.BlockId%>_probe_ccp_cachefill_doneId_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cachefill_done_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cache_evict_vld_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPDATA-1:0]         <%=obj.BlockId%>_probe_ccp_cache_evict_data_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPBYTEEN-1:0]       <%=obj.BlockId%>_probe_ccp_cache_evict_byten_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cache_evict_last_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cache_evict_cancel_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cache_evict_rdy_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cache_rdrsp_vld_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPDATA-1:0]         <%=obj.BlockId%>_probe_ccp_cache_rdrsp_data_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPBYTEEN-1:0]       <%=obj.BlockId%>_probe_ccp_cache_rdrsp_byten_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cache_rdrsp_last_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cache_rdrsp_cancel_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cache_rdrsp_rdy_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPADDR-1:0]         <%=obj.BlockId%>_probe_ccp_ctrlop_addr_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPSECURITY-1:0]     <%=obj.BlockId%>_probe_ccp_ctrlop_security_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPBANKBIT-1:0]      <%=obj.BlockId%>_probe_ccp_ctrlop_rdy_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_ctrlop_allocate_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_ctrlop_rd_data_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_ctrlop_wr_data_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_ctrlop_port_sel_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_ctrlop_bypass_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_ctrlop_rp_update_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_ctrlop_cancel_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_ctrlop_tag_state_update_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPBUSRTLN-1:0]      <%=obj.BlockId%>_probe_ccp_ctrlop_burstln_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_ctrlop_burstwrap_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_ctrlop_setway_debug_t;
typedef bit [<%=obj.nWays%>-1:0]            <%=obj.BlockId%>_probe_ccp_ctrlop_waybusy_vec_t;
typedef bit [<%=obj.nWays%>-1:0]            <%=obj.BlockId%>_probe_ccp_ctrlop_waystale_vec_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPBANKBIT-1:0]      <%=obj.BlockId%>_probe_ccp_cacheop_rdy_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cache_vld_t;
typedef bit [<%=obj.nWays%>-1:0]            <%=obj.BlockId%>_probe_ccp_cache_alloc_wayn_t;
typedef bit [<%=obj.nWays%>-1:0]            <%=obj.BlockId%>_probe_ccp_cache_hit_wayn_t;
typedef bit [<%=obj.nWays%>-1:0]            <%=obj.BlockId%>_probe_ccp_cache_wayn_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cache_evictvld_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPADDR-1:0]         <%=obj.BlockId%>_probe_ccp_cache_evictaddr_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPSECURITY-1:0]     <%=obj.BlockId%>_probe_ccp_cache_evictsecurity_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cache_nackuce_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cache_nack_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cache_nackce_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cachenacknoalloc_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_cachenoways2alloc_t;
//scratchpad related data types
typedef logic [<%=obj.nDataBanks%>-1:0]                        <%=obj.BlockId%>_probe_ccp_sp_ctrl_rdy_logic_t;  
typedef logic [<%=obj.nDataBanks%>-1:0]                        <%=obj.BlockId%>_probe_ccp_sp_ctrl_vld_logic_t ;      
typedef logic                                                  <%=obj.BlockId%>_probe_ccp_sp_ctrl_wr_data_logic_t;
typedef logic                                                  <%=obj.BlockId%>_probe_ccp_sp_ctrl_rd_data_logic_t;  
typedef logic [$clog2(<%=obj.nSets%>/<%=obj.nDataBanks%>)-1:0] <%=obj.BlockId%>_probe_ccp_sp_ctrl_index_addr_logic_t;
typedef logic [$clog2(<%=obj.nDataBanks%>)-1:0]                <%=obj.BlockId%>_probe_ccp_sp_ctrl_data_bank_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPWAYS-1:0]                                   <%=obj.BlockId%>_probe_ccp_sp_ctrl_way_num_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPBEAT-1:0]                                   <%=obj.BlockId%>_probe_ccp_sp_ctrl_beat_num_logic_t; 
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPBUSRTLN-1:0]                                <%=obj.BlockId%>_probe_ccp_sp_ctrl_burst_len_logic_t;
typedef logic                                                  <%=obj.BlockId%>_probe_ccp_sp_ctrl_burst_type_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WSMIMSG-1:0]                                    <%=obj.BlockId%>_probe_ccp_sp_ctrl_msg_type_logic_t;
typedef bit [<%=obj.nDataBanks%>-1:0]                        <%=obj.BlockId%>_probe_ccp_sp_ctrl_rdy_t;
typedef bit [<%=obj.nDataBanks%>-1:0]                        <%=obj.BlockId%>_probe_ccp_sp_ctrl_vld_t;      
typedef bit                                                  <%=obj.BlockId%>_probe_ccp_sp_ctrl_wr_data_t;
typedef bit                                                  <%=obj.BlockId%>_probe_ccp_sp_ctrl_rd_data_t;  
typedef bit [$clog2(<%=obj.nSets%>/<%=obj.nDataBanks%>)-1:0] <%=obj.BlockId%>_probe_ccp_sp_ctrl_index_addr_t;
typedef bit [$clog2(<%=obj.nDataBanks%>)-1:0]                <%=obj.BlockId%>_probe_ccp_sp_ctrl_data_bank_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPWAYS-1:0]                                   <%=obj.BlockId%>_probe_ccp_sp_ctrl_way_num_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPBEAT-1:0]                                   <%=obj.BlockId%>_probe_ccp_sp_ctrl_beat_num_t; 
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPBUSRTLN-1:0]                                <%=obj.BlockId%>_probe_ccp_sp_ctrl_burst_len_t;
typedef bit                                                  <%=obj.BlockId%>_probe_ccp_sp_ctrl_burst_type_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WSMIMSG-1:0]                                    <%=obj.BlockId%>_probe_ccp_sp_ctrl_msg_type_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCSRDATA-1:0]         <%=obj.BlockId%>_probe_ccp_csr_maint_wrdata_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCSRDATA-1:0]         <%=obj.BlockId%>_probe_ccp_csr_maint_rddata_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCSRDATA-1:0]         <%=obj.BlockId%>_probe_ccp_csr_maint_req_data_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCSROP-1:0]           <%=obj.BlockId%>_probe_ccp_csr_maint_req_opc_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCSRWAY-1:0]          <%=obj.BlockId%>_probe_ccp_csr_maint_req_way_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCSRENTRY-1:0]        <%=obj.BlockId%>_probe_ccp_csr_maint_req_entry_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCSRWORD-1:0]         <%=obj.BlockId%>_probe_ccp_csr_maint_req_word_t;
typedef bit [<%=obj.BlockId%>_probe_ccp_WCCPARRAYSEL-1:0]     <%=obj.BlockId%>_probe_ccp_csr_maint_req_array_sel_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_csr_maint_active_t;
typedef bit                        <%=obj.BlockId%>_probe_ccp_csr_maint_rddata_en_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPDATA_IF-1:0]      <%=obj.BlockId%>_probe_ccp_ctrlwr_data_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_ctrlwr_vld_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPBYTEEN-1:0]       <%=obj.BlockId%>_probe_ccp_ctrlwr_byten_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPBEAT-1:0]         <%=obj.BlockId%>_probe_ccp_ctrlwr_beatn_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_ctrlwr_last_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cachewr_rdy_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_ctrlfilldata_vld_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPDATA_IF-1:0]      <%=obj.BlockId%>_probe_ccp_ctrlfill_data_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPFILLID-1:0]       <%=obj.BlockId%>_probe_ccp_ctrlfilldata_Id_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPADDR-1:0]         <%=obj.BlockId%>_probe_ccp_ctrlfilldata_addr_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPWAYS-1:0]         <%=obj.BlockId%>_probe_ccp_ctrlfilldata_wayn_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPBEAT-1:0]         <%=obj.BlockId%>_probe_ccp_ctrlfilldata_beatn_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPBYTEEN-1:0]       <%=obj.BlockId%>_probe_ccp_ctrlfilldata_byten_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_ctrlfilldata_last_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cachefilldata_rdy_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_ctrlfill_vld_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPADDR-1:0]         <%=obj.BlockId%>_probe_ccp_ctrlfill_addr_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPWAYS-1:0]         <%=obj.BlockId%>_probe_ccp_ctrlfill_wayn_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPSECURITY-1:0]     <%=obj.BlockId%>_probe_ccp_ctrlfill_security_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPCACHESTATE-1:0]   <%=obj.BlockId%>_probe_ccp_ctrlfill_state_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cachefill_rdy_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPFILLDONEID-1:0]   <%=obj.BlockId%>_probe_ccp_cachefill_doneId_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cachefill_done_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cache_evict_vld_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPDATA_IF-1:0]      <%=obj.BlockId%>_probe_ccp_cache_evict_data_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPBYTEEN-1:0]       <%=obj.BlockId%>_probe_ccp_cache_evict_byten_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cache_evict_last_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cache_evict_cancel_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cache_evict_rdy_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cache_rdrsp_vld_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPDATA_IF-1:0]      <%=obj.BlockId%>_probe_ccp_cache_rdrsp_data_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPBYTEEN-1:0]       <%=obj.BlockId%>_probe_ccp_cache_rdrsp_byten_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cache_rdrsp_last_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cache_rdrsp_cancel_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cache_rdrsp_rdy_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPBANKBIT-1:0]      <%=obj.BlockId%>_probe_ccp_ctrlop_vld_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPADDR-1:0]         <%=obj.BlockId%>_probe_ccp_ctrlop_addr_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPSECURITY-1:0]     <%=obj.BlockId%>_probe_ccp_ctrlop_security_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPBANKBIT-1:0]      <%=obj.BlockId%>_probe_ccp_ctrlop_rdy_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_ctrlop_allocate_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_ctrlop_rd_data_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_ctrlop_wr_data_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_ctrlop_port_sel_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_ctrlop_bypass_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_ctrlop_rp_update_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_ctrlop_tagstateup_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPBUSRTLN-1:0]      <%=obj.BlockId%>_probe_ccp_ctrlop_burstln_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_ctrlop_burstwrap_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_ctrlop_setway_debug_logic_t;
typedef logic [<%=obj.nWays%>-1:0]            <%=obj.BlockId%>_probe_ccp_ctrlop_waybusy_vec_logic_t;
typedef logic [<%=obj.nWays%>-1:0]            <%=obj.BlockId%>_probe_ccp_ctrlop_waystale_vec_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPBANKBIT-1:0]      <%=obj.BlockId%>_probe_ccp_cacheop_rdy_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cache_vld_logic_t;
typedef logic [<%=obj.nWays%>-1:0]            <%=obj.BlockId%>_probe_ccp_cache_alloc_wayn_logic_t;
typedef logic [<%=obj.nWays%>-1:0]            <%=obj.BlockId%>_probe_ccp_cache_hit_wayn_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cache_evictvld_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPADDR-1:0]         <%=obj.BlockId%>_probe_ccp_cache_evictaddr_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cache_nackuce_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cache_nack_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cache_nackce_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cachenacknoalloc_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_cachenoways2alloc_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCSRDATA-1:0]        <%=obj.BlockId%>_probe_ccp_csr_maint_wrdata_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCSRDATA-1:0]        <%=obj.BlockId%>_probe_ccp_csr_maint_req_data_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCSRDATA-1:0]        <%=obj.BlockId%>_probe_ccp_csr_maint_rddata_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCSROP-1:0]          <%=obj.BlockId%>_probe_ccp_csr_maint_req_opc_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCSRWAY-1:0]         <%=obj.BlockId%>_probe_ccp_csr_maint_req_way_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCSRENTRY-1:0]       <%=obj.BlockId%>_probe_ccp_csr_maint_req_entry_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCSRWORD-1:0]        <%=obj.BlockId%>_probe_ccp_csr_maint_req_word_logic_t;
typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPARRAYSEL-1:0]    <%=obj.BlockId%>_probe_ccp_csr_maint_req_array_sel_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_csr_maint_active_logic_t;
typedef logic                        <%=obj.BlockId%>_probe_ccp_csr_maint_rddata_en_logic_t;

typedef logic [<%=obj.BlockId%>_probe_ccp_WCCPCACHESTATE-1:0]   <%=obj.BlockId%>_probe_ccp_cachestate_logic_t; 

/*
 <%=JSON.stringify(obj,null,' ')%>
 */

<% } %>
