`include "chi_coh_entry_virtual_seq.sv"
`include "chi_linkup_virtual_seq.sv"
`include "chi_coh_bringup_virtual_seq.sv"
