`ifdef USE_VIP_SNPS

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import svt_uvm_pkg::*;
  // Import the AMBA VIP
  import svt_amba_uvm_pkg::*;
`endif // USE_VIP_SNPS
