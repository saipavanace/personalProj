
//FileName: concerto_system_pkg.sv
//FIXME: Temp package
package concerto_system_pkg;

`include "concerto_system_params.svh"
`include "concerto_system_phys.svh"

endpackage: concerto_system_pkg
