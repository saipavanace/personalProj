//`ifdef USE_VIP_SNPS

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import svt_uvm_pkg::*;
  //import svt_chi_uvm_pkg::*;
  import svt_amba_uvm_pkg::*;
  /** Import the AMBA COMMON Package for amba_pv_extension */
  //import svt_amba_common_uvm_pkg::*;

//`endif // USE_VIP_SNPS
