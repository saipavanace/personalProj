////////////////////////////
//Description: Inlucde all AIU tests in this file
//File: aiu_test_lib.svh
////////////////////////////
`include "base_test.sv"
`include "bring_up_test.sv"
`include "ioaiu_qchannel_test.sv"
