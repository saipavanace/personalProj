// Library of all virtual sequences used in CHI Subsystem
`include "chi_subsys_base_vseq.sv"
`include "chi_subsys_dvmop_vseq.sv"
`include "chi_subsys_mkrdunq_error_vseq.sv"
`include "chi_subsys_write_excl_vseq.sv"
`include "chi_subsys_excl_noncoh_fix_addr_vseq.sv"
`include "chi_subsys_comb_wrcmo_vseq.sv"
`include "chi_subsys_unsupported_txn_vseq.sv"
`include "chi_subsys_atomic_stress_vseq.sv"
`include "chi_subsys_stash_stress_vseq.sv"
`include "chi_subsys_ip_error_vseq.sv"
`include "chi_subsys_random_vseq.sv"
`include "chi_subsys_random_native_interface_delay_vseq.sv"
`include "chi_subsys_error_vseq.sv"
`include "chi_subsys_snp_vseq.sv"
`include "chi_subsys_perf_vseq.sv"
`include "chi_subsys_random_noncoh_vseq.sv"
`include "chi_subsys_random_coherency_vseq.sv"
`include "chi_subsys_directed_noncoh_wr_rd_check_vseq.sv"
`include "chi_subsys_multicopy_atomicity_check_vseq.sv"
`include "chi_subsys_directed_atomic_self_check_vseq.sv"
`include "chi_subsys_directed_coh_wr_rd_check_vseq.sv"
`include "chi_subsys_cmo_vseq.sv"
`include "chi_subsys_mkrdunq_vseq.sv"
`include "chi_subsys_wrevctorevct_vseq.sv"
`include "chi_subsys_directed_atomic_vseq.sv"
`include "chi_subsys_vseq.sv" // USE in CASE of EMULATION
