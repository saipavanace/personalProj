//////////////////////////TB_  IRQ_if ////////////////////////
//DUT interfaces
//////////////////////////////////////////////////////////////////
interface IRQ_if;

  wire IRQ_c; 
  wire IRQ_uc;
  
endinterface: IRQ_if

