////////////////////////////////////////////////////////////////////////////////
//
// Cache State Test Generator Package
//
////////////////////////////////////////////////////////////////////////////////

package <%=obj.BlockId%>_CacheStateTestGenPkg;

import <%=obj.BlockId%>_ConcertoPkg::*;

`include "<%=obj.BlockId%>_CacheStateTestGen.svh"
`include "<%=obj.BlockId%>_AceStateTestGen.svh"

endpackage : <%=obj.BlockId%>_CacheStateTestGenPkg
