`timescale 1 ns/1 ps

<% if(obj.useResiliency) { %>
`include "fault_injector_checker.sv"
`include "placeholder_connectivity_checker.sv"
<% } %>
`ifdef USE_VIP_SNPS
   `include "snps_compile.sv"  
    `include "<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_connect_source2target_if.sv"
    import wrapper_pkg_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>::*;
`endif
`ifdef USE_VIP_SNPS_APB
	`include "<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_connection_wrapper_to_svt_apb_if.sv"
`endif

 <%
     var useAceQosPort    = obj.DiiInfo[obj.Id].interfaces.axiInt.params.useQosPort;
     var useAceRegionPort = obj.DiiInfo[obj.Id].interfaces.axiInt.params.useRegionPort;
     var useAceCache      = obj.DiiInfo[obj.Id].interfaces.axiInt.params.useAceCache     ;
     var useAceProt       = obj.DiiInfo[obj.Id].interfaces.axiInt.params.useProtPort     ;
     var useAceQos        = obj.DiiInfo[obj.Id].interfaces.axiInt.params.useQosPort      ;
     var useAceRegion     = obj.DiiInfo[obj.Id].interfaces.axiInt.params.useRegionPort   ;
     var useAceDomain     = obj.DiiInfo[obj.Id].interfaces.axiInt.params.useDomainPort   ;
     var wAwUser          = obj.DiiInfo[obj.Id].interfaces.axiInt.params.wAwUser    ;
     var wArUser          = obj.DiiInfo[obj.Id].interfaces.axiInt.params.wArUser    ;
     var wWUser           = obj.DiiInfo[obj.Id].interfaces.axiInt.params.wWUser     ;
     var wBUser           = obj.DiiInfo[obj.Id].interfaces.axiInt.params.wBUser     ;
     var wRUser           = obj.DiiInfo[obj.Id].interfaces.axiInt.params.wRUser     ;
   %>
module tb_top;


//-----------------------------------------------------------------------------
// Test and Env packages
//-----------------------------------------------------------------------------
import uvm_pkg::*;
<% if(obj.testBench == 'dii') { %>
`ifdef CDNS
`include "cdnAxiUvmDefines.sv"
import cdns_assert2uvm_pkg::*;
import DenaliSvCdn_axi::*;
import CdnSvVip::*;
import DenaliSvMem::*;
import DenaliSvChi::*;
import cdnChiUvm::*;
import cdnAxiUvm::*;
`endif // `ifndef CDNS
<% }  %>

import <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_test_lib_pkg::*;
import <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_env_pkg::*;

import <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_smi_agent_pkg::*;   //to get the *_FUNIT_IDS 
`include "snps_import.sv"
//-----------------------------------------------------------------------------
// vars
//-----------------------------------------------------------------------------

// Clocks and Reset
logic dut_clk;
logic tb_clk;
logic fr_clk;
logic tb_rstn;
logic temp_tb_rstn;
logic test_en;
logic soft_rstn;
logic reset_n_1d;



//error
int singleBitPct, doubleBitPct;

<% if(obj.useResiliency) { %>
 logic[1023:0] slv_req_corruption_vector = 1024'b0;
 logic[1023:0] slv_data_corruption_vector = 1024'b0;
 logic[WSMIADDR-1:0] smi_req_addr_modified;
 logic[<%=obj.DiiInfo[obj.Id].wData%>-1:0] smi_req_data_modified;  //TODO checkme: flat view of txn payload data for error injection

 logic bist_bist_next;
 logic bist_bist_next_ack;
 logic bist_domain_is_on;
 logic fault_mission_fault;
 logic fault_latent_fault;
 logic fault_cerr_over_thres_fault;
<% } %>

// Pipelined signals
logic CECR_ErrDetEn_1d;
logic UECR_ErrDetEn_1d;

//----------------------------------------------------------------------------
// Interfaces
//----------------------------------------------------------------------------
<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_stall_if <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if(); // PERF_CNT STALL_IF
initial uvm_config_db#(virtual <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_stall_if)::set(null, "", "<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_m_top_stall_if",       <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if); 

// Latency if
<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_latency_if <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_latency_if(); // PERF_CNT Latency_IF
initial uvm_config_db#(virtual <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_latency_if)::set(null, "", "<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_m_top_latency_if",       <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_latency_if); 

<%for(var i = 0; i < obj.DiiInfo[obj.Id].interfaces.smiTxInt.length; i++) { %>
<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_smi_if  m_smi<%=i%>_rx_smi_if(dut_clk, soft_rstn, "m_smi<%=i%>_rx_smi_if");
<% } %>
<%for(var i = 0; i < obj.DiiInfo[obj.Id].interfaces.smiRxInt.length; i++) { %>
<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_smi_if  m_smi<%=i%>_tx_smi_if(dut_clk, soft_rstn, "m_smi<%=i%>_tx_smi_if");
<% } %>

//`ifdef INHOUSE_AXI
<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_if m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if(dut_clk, soft_rstn);
<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_apb_if     m_apb_if(dut_clk, soft_rstn);
//`else
// SNPS AXI VIP inteface
`ifdef USE_VIP_SNPS
svt_axi_if axi_vip_if();

assign axi_vip_if.slave_if[0].aresetn = soft_rstn;
assign axi_vip_if.common_aclk = dut_clk;

<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_connect_source2target_slv_if m_wrapper_axi_inst (m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if, axi_vip_if.slave_if[0]);
`endif //  `ifdef USE_VIP_SNPS
`ifdef USE_VIP_SNPS_APB
svt_apb_if apb_vip_if();
assign apb_vip_if.pclk = dut_clk;
assign apb_vip_if.presetn = soft_rstn;
<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_connection_wrapper_to_svt_apb_if m_wrapper_apb_inst(m_apb_if,apb_vip_if);
`endif

<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_dii_rtl_if m_dii_rtl_if(dut_clk, soft_rstn);


//Q-channel interface
<%=obj.BlockId%>_q_chnl_if  m_q_chnl_if(fr_clk, tb_rstn);

uvm_event         toggle_clk;
uvm_event         toggle_rstn;
uvm_event         system_quiesce;
uvm_event         system_unquiesce;

uvm_event         injectSingleErrRtt;
uvm_event         injectDoubleErrRtt;

uvm_event         checkCELR;
uvm_event         checkUELR;

uvm_event         forceClkgate;
uvm_event         releaseClkgate;;

initial begin
   toggle_clk = new("toggle_clk");
   uvm_config_db#(uvm_event)::set(.cntxt( uvm_root::get()),
                                  .inst_name( "" ),
                                  .field_name( "toggle_clk" ),
                                  .value(toggle_clk));
   toggle_rstn = new("toggle_rstn");
   uvm_config_db#(uvm_event)::set(.cntxt( uvm_root::get()),
                                  .inst_name( "" ),
                                  .field_name( "toggle_rstn" ),
                                  .value(toggle_rstn));
end

bit enable=1;
always @(posedge fr_clk) begin
    toggle_clk.wait_trigger();
    @(negedge fr_clk);
    $display("triggered toggle_clk_event @time: %0t",$time);
    enable = ~enable;
end

assign dut_clk = enable ? fr_clk : 0;

bit soft_rstn_en=1;
always @(posedge fr_clk) begin
    toggle_rstn.wait_trigger();
    @(negedge fr_clk);
    $display("treggered reset event @time: %0t",$time);
    soft_rstn_en = ~soft_rstn_en;
end

// delay tb_rstn to allow test_en to toggle
initial begin
   test_en = 1'b1;
   tb_rstn = 1'b0;
end

always @(posedge temp_tb_rstn) begin
   test_en = 1'b0;
   repeat (5) @(negedge fr_clk);
   tb_rstn = ~tb_rstn;
end

assign soft_rstn = soft_rstn_en ? tb_rstn : 0;

`ifdef RTL_DUT

//--------------------------------------------------------------------------
//instantiate and connect dut
//--------------------------------------------------------------------------

<% if(obj.useResiliency) { %>
assign bist_bist_next = 1'b0;
<% } %>
<% if ( obj.DiiInfo[obj.Id].configuration ) { %>
config_dii_a dut
<% } else if(obj.instanceName) { %>
<%=obj.instanceMap[obj.instanceName]%> dut
<% } else { %>						      
dii_top_0 dut
<% } %>  
     (
    //HW layer signals **********************************************************
    .<%=obj.DiiInfo[obj.Id].interfaces.clkInt.name%>clk(dut_clk),

    .<%=obj.DiiInfo[obj.Id].interfaces.uIdInt.name%>my_f_unit_id(<%=obj.DiiInfo[obj.Id].interfaces.uIdInt.params.wFUnitId%>'d<%=obj.DiiInfo[obj.Id].FUnitId%>),   //from js config
    .<%=obj.DiiInfo[obj.Id].interfaces.uIdInt.name%>my_n_unit_id(<%=obj.DiiInfo[obj.Id].interfaces.uIdInt.params.wNUnitId%>'d<%=obj.DiiInfo[obj.Id].nUnitId%>),   //from js config
    .<%=obj.DiiInfo[obj.Id].interfaces.uIdInt.name%>my_csr_rpn(<%=obj.DiiInfo[obj.Id].interfaces.uIdInt.params.wRpn%>'d<%=obj.DiiInfo[obj.Id].rpn%>),             //from js config
    .<%=obj.DiiInfo[obj.Id].interfaces.uIdInt.name%>my_csr_nrri(<%=obj.DiiInfo[obj.Id].interfaces.uIdInt.params.wNrri%>'d<%=obj.DiiInfo[obj.Id].nrri%>),          //from js config
      
<% if(obj.useResiliency) { %>
    //TODO resiliency if ******************************************
<% if(obj.DiiInfo[obj.Id].ResilienceInfo.enableUnitDuplication) { %>
    .<%=obj.DiiInfo[obj.Id].interfaces.checkClkInt.name%>clk(dut_clk),
    .<%=obj.DiiInfo[obj.Id].interfaces.checkClkInt.name%>test_en(test_en),
//    .<%=obj.DiiInfo[obj.Id].interfaces.checkClkInt.name%>reset_n(soft_rstn),
<% } %>
<% if (!obj.DiiInfo[obj.Id].interfaces.bistDebugDisableInt._SKIP_) { %>
    .<%=obj.DiiInfo[obj.Id].interfaces.bistDebugDisableInt.name%>pin     ('h1),
<% } %>
    // .clk_check(fr_clk),
     .bist_bist_next(bist_bist_next),
     .bist_bist_next_ack(bist_bist_next_ack),
     .bist_domain_is_on(bist_domain_is_on),
     .fault_mission_fault(fault_mission_fault),
     .fault_latent_fault(fault_latent_fault),
     .fault_cerr_over_thres_fault(fault_cerr_over_thres_fault),
<% } %>

    //APB control if *****************************************
    .<%=obj.DiiInfo[obj.Id].interfaces.apbInt.name%>paddr        (m_apb_if.paddr[<%=obj.DiiInfo[obj.Id].interfaces.apbInt.params.wAddr%>-1:0]),
    .<%=obj.DiiInfo[obj.Id].interfaces.apbInt.name%>pwrite       (m_apb_if.pwrite),
    .<%=obj.DiiInfo[obj.Id].interfaces.apbInt.name%>psel         (m_apb_if.psel),
    .<%=obj.DiiInfo[obj.Id].interfaces.apbInt.name%>penable      (m_apb_if.penable),
    .<%=obj.DiiInfo[obj.Id].interfaces.apbInt.name%>prdata       (m_apb_if.prdata),
    .<%=obj.DiiInfo[obj.Id].interfaces.apbInt.name%>pwdata       (m_apb_if.pwdata),
    .<%=obj.DiiInfo[obj.Id].interfaces.apbInt.name%>pready       (m_apb_if.pready),
    .<%=obj.DiiInfo[obj.Id].interfaces.apbInt.name%>pslverr      (m_apb_if.pslverr),
<%  if(obj.DiiInfo[obj.Id].interfaces.apbInt.params.wProt !== 0) { %>
    .<%=obj.DiiInfo[obj.Id].interfaces.apbInt.name%>pprot        (m_apb_if.pprot),
<% } %>
<%  if(obj.DiiInfo[obj.Id].interfaces.apbInt.params.wStrb !== 0) { %>
    .<%=obj.DiiInfo[obj.Id].interfaces.apbInt.name%>pstrb        (m_apb_if.pstrb),
<% } %>
    .<%=obj.DiiInfo[obj.Id].interfaces.irqInt.name%>c            (m_apb_if.IRQ_c),
    .<%=obj.DiiInfo[obj.Id].interfaces.irqInt.name%>uc           (m_apb_if.IRQ_uc),



    //SMI ***************************************************

<%for (var i = 0; i < obj.DiiInfo[obj.Id].interfaces.smiTxInt.length; i++) { %>
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>ndp_msg_valid         (m_smi<%=i%>_rx_smi_if.smi_msg_valid ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>ndp_msg_ready         (m_smi<%=i%>_rx_smi_if.smi_msg_ready  ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>ndp_ndp_len           (m_smi<%=i%>_rx_smi_if.smi_ndp_len   ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>ndp_dp_present        (m_smi<%=i%>_rx_smi_if.smi_dp_present) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>ndp_targ_id           (m_smi<%=i%>_rx_smi_if.smi_targ_id   ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>ndp_src_id            (m_smi<%=i%>_rx_smi_if.smi_src_id    ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>ndp_msg_id            (m_smi<%=i%>_rx_smi_if.smi_msg_id    ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>ndp_msg_type          (m_smi<%=i%>_rx_smi_if.smi_msg_type  ) ,
<% if(obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].params.wSmiUser >0) {%>
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name %>ndp_msg_user         (m_smi<%=i%>_rx_smi_if.smi_msg_user  ) ,
<% } %>
<% if(obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].params.wSmiTier >0) {%>
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>ndp_msg_tier          (m_smi<%=i%>_rx_smi_if.smi_msg_tier  ) ,
<% } %>
<% if(obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].params.wSmiSteer >0) {%>
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>ndp_steer             (m_smi<%=i%>_rx_smi_if.smi_steer     ) ,
<% } %>
<% if(obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].params.wSmiPri >0) {%>
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>ndp_msg_pri           (m_smi<%=i%>_rx_smi_if.smi_msg_pri   ) ,
<% } %>
<% if(obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].params.wSmiMsgQos >0) {%>
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>ndp_msg_qos           (m_smi<%=i%>_rx_smi_if.smi_msg_qos   ) ,
<% } %>
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>ndp_ndp               (m_smi<%=i%>_rx_smi_if.smi_ndp[<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].params.wSmiNDP%>-1:0]) ,
<% if(obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].params.wSmiErr >0) {%>
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>ndp_msg_err           (m_smi<%=i%>_rx_smi_if.smi_msg_err   ) ,
<% } %>

 <%  if (obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].params.wSmiDPdata >0) { %>    
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>dp_valid              (m_smi<%=i%>_rx_smi_if.smi_dp_valid  ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>dp_ready              (m_smi<%=i%>_rx_smi_if.smi_dp_ready  ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>dp_last               (m_smi<%=i%>_rx_smi_if.smi_dp_last   ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>dp_data               (m_smi<%=i%>_rx_smi_if.smi_dp_data   ) ,
<% if(obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].params.wSmiDPuser >0) {%>
.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>dp_user               (m_smi<%=i%>_rx_smi_if.smi_dp_user   ) ,
<% } %>

    <% } %>
<% } %>
<%for (var i = 0; i < obj.DiiInfo[obj.Id].interfaces.smiRxInt.length; i++) { %>
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_msg_valid         (m_smi<%=i%>_tx_smi_if.smi_msg_valid ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_msg_ready         (m_smi<%=i%>_tx_smi_if.smi_msg_ready ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_ndp_len           (m_smi<%=i%>_tx_smi_if.smi_ndp_len   ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_dp_present        (m_smi<%=i%>_tx_smi_if.smi_dp_present) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_targ_id           (m_smi<%=i%>_tx_smi_if.smi_targ_id   ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_src_id            (m_smi<%=i%>_tx_smi_if.smi_src_id    ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_msg_id            (m_smi<%=i%>_tx_smi_if.smi_msg_id    ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_msg_type          (m_smi<%=i%>_tx_smi_if.smi_msg_type  ) ,
<% if(obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].params.wSmiUser >0) {%>
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_msg_user          (m_smi<%=i%>_tx_smi_if.smi_msg_user  ) ,
<% } %>
<% if(obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].params.wSmiTier >0) {%>
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_msg_tier          (m_smi<%=i%>_tx_smi_if.smi_msg_tier  ) ,
<% } %>
<% if(obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].params.wSmiSteer >0) {%>
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_steer             (m_smi<%=i%>_tx_smi_if.smi_steer     ) ,
<% } %>
<% if(obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].params.wSmiPri >0) {%>
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_msg_pri           (m_smi<%=i%>_tx_smi_if.smi_msg_pri   ) ,
<% } %>
<% if(obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].params.wSmiMsgQos >0) {%>
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_msg_qos           (m_smi<%=i%>_tx_smi_if.smi_msg_qos   ) ,
<% } %>
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_ndp               (m_smi<%=i%>_tx_smi_if.smi_ndp[<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].params.wSmiNDP%>-1:0]) ,
<% if(obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].params.wSmiErr >0) {%>
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_msg_err           (m_smi<%=i%>_tx_smi_if.smi_msg_err   ) ,
<% } %>
    <%  if (obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].params.wSmiDPdata >0) { %>    
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>dp_valid              (m_smi<%=i%>_tx_smi_if.smi_dp_valid  ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>dp_ready              (m_smi<%=i%>_tx_smi_if.smi_dp_ready  ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>dp_last               (m_smi<%=i%>_tx_smi_if.smi_dp_last   ) ,
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>dp_data               (m_smi<%=i%>_tx_smi_if.smi_dp_data   ) ,
<% if(obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].params.wSmiDPuser >0) {%>
.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>dp_user               (m_smi<%=i%>_tx_smi_if.smi_dp_user   ) ,
<% } %>
    <% } %>
<% } %>
    // Trace-Debug (DVE ID) ***********************************************
<% if(obj.testBench == 'dii') { %>
`ifdef CDNS
.<%=obj.DiiInfo[obj.Id].interfaces.uSysDveIdInt.name%>f_unit_id            ('{(<%=obj.DveInfo[0].interfaces.uIdInt.params.wFUnitId%>){<%=obj.DveInfo[0].FUnitId%>}} ),
`else
.<%=obj.DiiInfo[obj.Id].interfaces.uSysDveIdInt.name%>f_unit_id            ({(<%=obj.DveInfo[0].interfaces.uIdInt.params.wFUnitId%>){<%=obj.DveInfo[0].FUnitId%>}} ),
`endif // `ifndef CDNS
<% } else {%>
.<%=obj.DiiInfo[obj.Id].interfaces.uSysDveIdInt.name%>f_unit_id            ({(<%=obj.DveInfo[0].interfaces.uIdInt.params.wFUnitId%>){<%=obj.DveInfo[0].FUnitId%>}} ),
<% } %>
      
    // AXI ****************************************************************
 //`ifdef INHOUSE_AXI
<% if(obj.DiiInfo[obj.Id].interfaces.axiInt.params.wProt) { %>
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>aw_prot        ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awprot              ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>ar_prot        ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arprot              ) ,
<% } %>
<%if (obj.DiiInfo[obj.Id].interfaces.axiInt.params.wQos){%>
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>aw_qos         ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awqos               ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>ar_qos         ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arqos               ) ,
<% } %>
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>aw_ready       ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awready             ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>aw_valid       ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awvalid             ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>aw_id          ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awid  [<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wAwId%>-1:0]       ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>aw_addr        ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awaddr[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wAddr%>-1:0]       ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>aw_burst       ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awburst             ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>aw_len         ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awlen [<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wLen%> -1:0]       ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>aw_lock        ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awlock[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wLock%>-1:0]       ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>aw_size        ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awsize[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wSize%>-1:0]       ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>w_ready        ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.wready              ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>w_valid        ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.wvalid              ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>w_data         ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.wdata[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wData%>-1:0]        ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>w_last         ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.wlast               ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>w_strb         ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.wstrb[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wData%>/8-1:0]      ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>b_ready        ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.bready              ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>b_valid        ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.bvalid              ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>b_id           ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.bid  [<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wAwId%>-1:0]        ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>b_resp         ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.bresp[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wResp%>-1:0]        ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>ar_ready       ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arready             ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>ar_valid       ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arvalid             ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>ar_addr        ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.araddr[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wAddr%>-1:0]       ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>ar_burst       ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arburst             ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>ar_id          ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arid  [<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wArId%>-1:0]       ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>ar_len         ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arlen [<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wLen%> -1:0]       ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>ar_lock        ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arlock[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wLock%>-1:0]       ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>ar_size        ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arsize[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wSize%>-1:0]       ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>r_id           ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.rid                 ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>r_resp         ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.rresp[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wResp%> -1:0]       ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>r_ready        ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.rready              ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>r_valid        ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.rvalid              ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>r_data         ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.rdata[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wData%> -1:0]       ) ,
     .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>r_last         ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.rlast               ) ,
    .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>aw_cache        ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awcache             ) ,
    .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>ar_cache        ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arcache             ) ,
<%if (obj.DiiInfo[obj.Id].interfaces.axiInt.wRegion){%>
    .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>aw_region       ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awregion[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wRegion%>-1:0]    ) ,
    .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>ar_region       ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arregion[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wRegion%>-1:0]    ) ,
<% } %>
<%if (wAwUser >0){%>
    .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>aw_user         ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awuser  [<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wAwUser%>-1:0]    ) ,
<% } %>
<%if (wWUser >0){%>
    .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>w_user          ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.wuser[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wWUser%>    -1:0]    ) ,
<% } %>
<%if (wBUser){%>
    .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>b_user          ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.buser[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wBUser%>    -1:0]    ) ,
<% } %>
<%if (wArUser){%>
    .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>ar_user         ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.aruser[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wArUser%>  -1:0]    ) ,
<% } %>
<%if (wRUser){%>
    .<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>r_user          ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.ruser[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wArUser%>   -1:0]    ) ,
<% } %>
<%if (useAceDomain){%>
<% } %>
//Q-channel interface connection
<% if(obj.DiiInfo[obj.Id].usePma) { %>
    .<%=obj.DiiInfo[obj.Id].interfaces.qInt.name%>ACTIVE                ( m_q_chnl_if.QACTIVE ) ,
    .<%=obj.DiiInfo[obj.Id].interfaces.qInt.name%>DENY                  ( m_q_chnl_if.QDENY   ) ,
    .<%=obj.DiiInfo[obj.Id].interfaces.qInt.name%>REQn                  ( m_q_chnl_if.QREQn   ) ,
    .<%=obj.DiiInfo[obj.Id].interfaces.qInt.name%>ACCEPTn               ( m_q_chnl_if.QACCEPTn) ,
<% } %>
     // PERF MON MASTER ENABLE
    .trigger_trigger(<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.master_cnt_enable),
    
    .<%=obj.DiiInfo[obj.Id].interfaces.clkInt.name%>test_en(test_en),
    .<%=obj.DiiInfo[obj.Id].interfaces.clkInt.name%>reset_n(soft_rstn)
      );
`endif //  `ifdef RTL_DUT
<%if( obj.DiiInfo[obj.Id].nPerfCounters> 0) { %> 
/////////////////////// PERF_CNT CONNECT DUT to LATENCY LATENCY_IF////////////////////////////////////////////////////
<%if( obj.DiiInfo[obj.Id].nLatencyCounters > 0) { %> 
assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_latency_if.clk              =   dut_clk;
assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_latency_if.rst_n            =   soft_rstn;
assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_latency_if.alloc_if         =   dut.u_dii_unit.u_ncr_pmon.latency_counter_in_alloc;
assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_latency_if.dealloc_if       =   dut.u_dii_unit.u_ncr_pmon.latency_counter_in_dealloc;
assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_latency_if.dut_latency_bins =   dut.u_dii_unit.u_ncr_pmon.latency_bins;
assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_latency_if.div_clk_rtl      =   dut.u_dii_unit.u_ncr_pmon.latency_counter_table.divevt_clk;
<% } %>
/////////////////////// PERF_CNT CONNECT STALL_IF TO DUT////////////////////////////////////////////////////

  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.clk = dut_clk;
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.rst_n = soft_rstn;
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.trace_capture_busy = dut.u_dii_unit.trace_capture_busy;

  // SMI TX
  <%for (var i = 0; i < obj.DiiInfo[obj.Id].interfaces.smiTxInt.length; i++) { %>
  <%  if (obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].params.wSmiDPdata >0) { %>  
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.smi_tx<%=i%>_valid = dut.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>dp_valid ;       
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.smi_tx<%=i%>_ready = dut.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>dp_ready  ; 
  <% } else { %>  
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.smi_tx<%=i%>_valid = dut.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>ndp_msg_valid ;       
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.smi_tx<%=i%>_ready = dut.<%=obj.DiiInfo[obj.Id].interfaces.smiTxInt[i].name%>ndp_msg_ready  ;      
  <% } %>
  <% } %> 
  // SMI RX
  <%for (var i = 0; i < obj.DiiInfo[obj.Id].interfaces.smiTxInt.length; i++) { %>
  <%  if (obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].params.wSmiDPdata >0) { %> 
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.smi_rx<%=i%>_valid = dut.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>dp_valid;
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.smi_rx<%=i%>_ready = dut.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>dp_ready;
  assign (supply0, supply1) dut.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>dp_valid = m_smi<%=i%>_tx_smi_if.force_smi_msg_valid;  
  assign (supply0, supply1) dut.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>dp_ready = m_smi<%=i%>_tx_smi_if.force_smi_msg_ready;
  <% } else { %> 
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.smi_rx<%=i%>_valid = dut.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_msg_valid;
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.smi_rx<%=i%>_ready = dut.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_msg_ready; 

  assign (supply0, supply1) dut.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_msg_valid = m_smi<%=i%>_tx_smi_if.force_smi_msg_valid;
  assign (supply0, supply1)  dut.<%=obj.DiiInfo[obj.Id].interfaces.smiRxInt[i].name%>ndp_msg_ready = m_smi<%=i%>_tx_smi_if.force_smi_msg_ready; 
  <% } %>
  <% } %>
  // AXI 
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.axi_aw_valid = dut.<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>aw_valid;
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.axi_aw_ready = dut.<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>aw_ready;
  
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.axi_w_valid = dut.<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>w_valid;
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.axi_w_ready = dut.<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>w_ready;
  
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.axi_ar_valid = dut.<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>ar_valid;
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.axi_ar_ready = dut.<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>ar_ready;
  
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.axi_r_valid = dut.<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>r_valid;
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.axi_r_ready = dut.<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>r_ready;
  
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.axi_b_valid = dut.<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>b_valid;
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.axi_b_ready = dut.<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>b_ready;
  /////////////////////////////////// DII BW events //////////////////////////////////////////////////
  //dtr_req event
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.dtr_req_valid = dut.u_dii_unit.dtr_req_valid;
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.dtr_req_ready = dut.u_dii_unit.dtr_req_ready;
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.dtr_req_funit_id_if = (dut.u_dii_unit.dtr_req_target_id >> WSMINCOREPORTID);
  <%if (wArUser > 0){%>
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.dtr_req_user_bits_if = dut.u_dii_unit.pmon_dtr_req_user_bits; //dut.u_dii_unit.dtr_req_aux;
  <% } %>
  //dtw_req event
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.dtw_req_valid = dut.u_dii_unit.dtw_req_valid;
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.dtw_req_ready = dut.u_dii_unit.dtw_req_ready;
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.dtw_req_funit_id_if = (dut.u_dii_unit.dtw_req_initiator_id >> WSMINCOREPORTID);
  <%if (wAwUser > 0){%>
  assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.dtw_req_user_bits_if = dut.u_dii_unit.pmon_dtw_req_user_bits; //dut.u_dii_unit.dtw_req_aux;
  <% } %>
  /////////////////// END PERF_CNT STALL_IF ////////////////////////////////////////////////////
<%for (var i = 0; i < obj.DutInfo.nPerfCounters; i++) { %>
assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.cnt_reg_capture[<%=i%>].cnt_v     =  dut.u_dii_unit.dii_csr.dii_csr_gen.DIICNTVR<%=i%>_CountVal_out ;  
assign <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_sb_stall_if.cnt_reg_capture[<%=i%>].cnt_v_str =  dut.u_dii_unit.dii_csr.dii_csr_gen.DIICNTSR<%=i%>_CountSatVal_out;      
<% } %>
`ifdef INHOUSE_AXI
/////FOCE READ DATA CHANNEL ET B RESPENSE CHANNEL FOR PERFMON////////////////////
assign (supply0, supply1) dut.<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>b_ready  = m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.force_bready;  
assign (supply0, supply1) dut.<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>b_valid  = m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.force_bvalid;
assign (supply0, supply1) dut.<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>r_ready  = m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.force_rready;  
assign (supply0, supply1) dut.<%=obj.DiiInfo[obj.Id].interfaces.axiInt.name%>r_valid  = m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.force_rvalid;
`endif //  `ifdef INHOUSE_AXI
initial begin
    if ($test$plusargs("forced_stall")) begin
        $assertoff(0,m_smi0_tx_smi_if);
        $assertoff(0,m_smi1_tx_smi_if);
        $assertoff(0,m_smi2_tx_smi_if);
    end
end

<% } %>
//--------------------------------------------------------------------------
//instantiate and connect coverage for standard interfaces
//--------------------------------------------------------------------------

// ARM AXI Assertions
`ifdef ASSERT_ON
`ifndef ASSERT_OFF  
<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_Axi4PC_ace #(.ADDR_WIDTH(<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wAddr%>),
	     .WID_WIDTH( <%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wAwId%>),
	     .RID_WIDTH( <%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wArId%>),
	     .AWUSER_WIDTH( <%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wAwUser%>),
	     .WUSER_WIDTH( <%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wWUser%>),
	     .BUSER_WIDTH( <%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wBUser%>),
	     .ARUSER_WIDTH( <%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wArUser%>),
	     .RUSER_WIDTH( <%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wRUser%>),
	     .DATA_WIDTH(<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wData%>))
   m_axi4_arm_sva     (
   // Global Signals
   .ACLK                     ( dut_clk                           ) ,
   .ARESETn                  ( soft_rstn                          ) ,

   // Write Address Channel
   .AWID                     ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awid  [<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wAwId%>-1:0]       ) ,
   .AWADDR                   ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awaddr[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wAddr%>-1:0]       ) ,
   .AWLEN                    ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awlen [<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wLen%> -1:0]       ) ,
   .AWSIZE                   ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awsize[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wSize%>-1:0]       ) ,
   .AWBURST                  ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awburst          ) ,
   .AWLOCK                   ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awlock[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wLock%>-1:0]       ) ,
   .AWCACHE                  ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awcache          ) ,
<% if ( obj.DiiInfo[obj.Id].interfaces.axiInt.params.wAwUser > 0 ) { %>
   .AWUSER                   ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awuser[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wAwUser%>-1:0]     ) ,
<% } %>
<% if(useAceProt) { %>
   .AWPROT                   ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awprot[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wProt%>-1:0]       ) ,
<% } else { %>
   .AWPROT                   (                                                                                                         ) ,
<% } %>
<% if(useAceQos) { %>
   .AWQOS                    ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awqos [<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wQos%> -1:0]       ) ,
<% } else { %>
   .AWQOS                    (                                                                                                         ) ,
<% } %>
<% if(useAceRegion) { %>
   .AWREGION                 ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awregion[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wRegion%>-1:0]   ) ,
<% } else { %>
   .AWREGION                 (                                                                                                         ) ,
<% } %>
   .AWVALID                  ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awvalid          ) ,
   .AWREADY                  ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.awready          ) ,

   // Write Channel
   .WDATA                    ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.wdata[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wData%>  -1:0]      ) ,
   .WSTRB                    ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.wstrb[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wData%>/8-1:0]      ) ,
<% if (obj.DiiInfo[obj.Id].interfaces.axiInt.params.wWUser ) { %>
   .WUSER                    ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.wuser[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wWUser%> -1:0]      ) ,
<% } %>
   .WLAST                    ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.wlast               ) ,
   .WVALID                   ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.wvalid              ) ,
   .WREADY                   ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.wready              ) ,

   // Write Response Channel
   .BID                      ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.bid  [<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wAwId%>  -1:0]      ) ,
   .BRESP                    ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.bresp[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wResp%>  -1:0]      ) ,
<% if ( obj.DiiInfo[obj.Id].interfaces.axiInt.params.wBUser ) { %>
   .BUSER                    ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.buser[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wBUser%> -1:0]      ) ,
<% } %>
   .BVALID                   ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.bvalid              ) ,
   .BREADY                   ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.bready              ) ,

   // Read Address Channel
   .ARID                     ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arid  [<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wArId%> -1:0]      ) ,
   .ARADDR                   ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.araddr[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wAddr%> -1:0]      ) ,
   .ARLEN                    ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arlen [<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wLen%>  -1:0]      ) ,
   .ARSIZE                   ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arsize[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wSize%> -1:0]      ) ,
   .ARBURST                  ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arburst             ) ,
   .ARLOCK                   ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arlock[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wLock%> -1:0]      ) ,
   .ARCACHE                  ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arcache             ) ,
<% if ( obj.DiiInfo[obj.Id].interfaces.axiInt.params.wArUser ) { %>
   .ARUSER                   ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.aruser[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wArUser%>-1:0]     ) ,
<% } %>
<% if(useAceProt) { %>
   .ARPROT                   ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arprot[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wProt%> -1:0]      ) ,
<% } else { %>
   .ARPROT                   (                                                                                                         ) ,
<% } %>
<% if(useAceQos) { %>
   .ARQOS                    ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arqos [<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wQos%>  -1:0]      ) ,
<% } else { %>
   .ARQOS                    (                                                                                                         ) ,		   
<% } %>
<% if(useAceRegion) { %>
   .ARREGION                 ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arregion[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wRegion%>-1:0]   ) ,
<% } else { %>
   .ARREGION                 (                                                                                                         ) ,
<% } %>
   .ARVALID                  ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arvalid             ) ,
   .ARREADY                  ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.arready             ) ,

   //  Read Channel
   .RID                      ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.rid  [<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wArId%>  -1:0]      ) ,
   .RLAST                    ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.rlast               ) ,
   .RDATA                    ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.rdata[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wData%>  -1:0]      ) ,
   .RRESP                    ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.rresp[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wResp%>  -1:0]      ) ,
<% if ( obj.DiiInfo[obj.Id].interfaces.axiInt.params.wRUser ) { %>
   .RUSER                    ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.ruser[<%=obj.DiiInfo[obj.Id].interfaces.axiInt.params.wArUser%>-1:0]      ) ,
<% } %>
   .RVALID                   ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.rvalid              ) ,
   .RREADY                   ( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.rready              ) ,

   // Low Power Interface
   .CACTIVE                  ( <%=obj.DiiInfo[obj.Id].interfaces.qInt.params.wActive%>'b1                                              ) ,
   .CSYSREQ                  ( 1'b1                              ) ,
   .CSYSACK                  ( 1'b1                              )
) ;
initial begin
    if ($test$plusargs("forced_stall")) begin
        $assertoff(0,m_axi4_arm_sva);
    end
end
`endif //ASSERT_OFF
`endif //ASSERT_ON

//-----------------------------------------------------------------------------
// Generate clocks and reset
//-----------------------------------------------------------------------------
clk_rst_gen #(.CLK_PERIOD(<%=obj.Clocks[0].params.period%>)) cr_gen (.clk_fr(fr_clk), .clk_tb(tb_clk), .rst(temp_tb_rstn));

//-----------------------------------------------------------------------------
// Connect RTL internal signals to if
//-----------------------------------------------------------------------------

// interface to tap internal csr signal
<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_dii_csr_probe_if u_csr_probe_if(.clk(dut_clk),.resetn(soft_rstn));

//TODO FIXME quiesce without ocp, sfi
`include "concerto_quiesce.sv"
initial begin
    if ($test$plusargs("inject_ttdebug")) begin
        quiesce_system();
        system_quiesce.trigger();
        `uvm_info("tb_top", "saw system quiesce",UVM_MEDIUM)
        system_unquiesce.wait_ptrigger();
        `uvm_info("tb_top", "saw end of debug injection",UVM_MEDIUM)
        unquiesce_system();
    end
end


<% if(obj.useResiliency) { %>
 fault_injector_checker fault_inj_check(dut_clk, soft_rstn);
 placeholder_connectivity_checker placeholder_connec_chk(dut_clk, soft_rstn);
 initial begin
<% if(obj.testBench == 'dii') { %>
`ifndef VCS

    uvm_config_db#(event)::set(.cntxt(null),
                               .inst_name( "*" ),
                               .field_name( "kill_test" ),
                               .value(placeholder_connec_chk.kill_test));

    uvm_config_db#(event)::set(.cntxt(null),
                               .inst_name( "*" ),
                               .field_name( "raise_obj_for_resiliency_test" ),
                               .value(fault_inj_check.raise_obj_for_resiliency_test));

    uvm_config_db#(event)::set(.cntxt(null),
                               .inst_name( "*" ),
                               .field_name( "drop_obj_for_resiliency_test" ),
                               .value(fault_inj_check.drop_obj_for_resiliency_test));
`else // `ifndef VCS
    placeholder_connec_chk.kill_test = new("kill_test");
    fault_inj_check.raise_obj_for_resiliency_test = new("raise_obj_for_resiliency_test");
    fault_inj_check.drop_obj_for_resiliency_test = new("drop_obj_for_resiliency_test");

    uvm_config_db#(uvm_event)::set(.cntxt(null),
                               .inst_name( "*" ),
                               .field_name( "kill_test" ),
                               .value(placeholder_connec_chk.kill_test));

    uvm_config_db#(uvm_event)::set(.cntxt(null),
                               .inst_name( "*" ),
                               .field_name( "raise_obj_for_resiliency_test" ),
                               .value(fault_inj_check.raise_obj_for_resiliency_test));

    uvm_config_db#(uvm_event)::set(.cntxt(null),
                               .inst_name( "*" ),
                               .field_name( "drop_obj_for_resiliency_test" ),
                               .value(fault_inj_check.drop_obj_for_resiliency_test));
`endif // `ifndef VCS ... `else ... 
<% } else {%>

    uvm_config_db#(event)::set(.cntxt(null),
                               .inst_name( "*" ),
                               .field_name( "kill_test" ),
                               .value(placeholder_connec_chk.kill_test));

    uvm_config_db#(event)::set(.cntxt(null),
                               .inst_name( "*" ),
                               .field_name( "raise_obj_for_resiliency_test" ),
                               .value(fault_inj_check.raise_obj_for_resiliency_test));

    uvm_config_db#(event)::set(.cntxt(null),
                               .inst_name( "*" ),
                               .field_name( "drop_obj_for_resiliency_test" ),
                               .value(fault_inj_check.drop_obj_for_resiliency_test));
<% } %>
 end

 ////TODO FIXME inject error in which IF?
 //assign smi_req_addr_modified = smi_if.smi_addr ^ slv_req_corruption_vector;
 //assign smi_req_data_modified = smi_if.smi_dp_data ^ slv_data_corruption_vector;
<% } %>


initial begin

    uvm_config_db#(virtual <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_dii_csr_probe_if)::set(.cntxt( uvm_root::get() ),
                                        .inst_name( "" ),
                                        .field_name( "u_csr_probe_if" ),
                                        .value( u_csr_probe_if ));

    <% for (i=0; i<obj.DiiInfo[obj.Id].interfaces.smiTxInt.length; i++) { %>
    uvm_config_db#(virtual <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_smi_if)::set(.cntxt( null ),
                                        .inst_name( "*" ),
                                        .field_name( "m_smi<%=i%>_rx_smi_if" ),
                                        .value( m_smi<%=i%>_rx_smi_if ));
    <% } %>
    <% for (i=0; i<obj.DiiInfo[obj.Id].interfaces.smiRxInt.length; i++) { %>
    uvm_config_db#(virtual <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_smi_if)::set(.cntxt( null ),
                                        .inst_name( "*" ),
                                        .field_name( "m_smi<%=i%>_tx_smi_if" ),
                                        .value( m_smi<%=i%>_tx_smi_if ));
    <% } %>

    `ifdef USE_VIP_SNPS
         m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.IS_ACTIVE = 0;
    `else // !`ifdef USE_VIP_SNPS
    
         m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if.IS_ACTIVE = 1;
    `endif // !`ifdef USE_VIP_SNPS
    uvm_config_db#(virtual <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_if)::set(.cntxt( uvm_root::get() ),
                                        .inst_name( "" ),
                                        .field_name( "m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if" ),
                                        .value( m_<%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_axi_slv_if ));


`ifdef USE_VIP_SNPS
            uvm_config_db#(svt_axi_vif)::set(uvm_root::get(), 
            "", "vif", axi_vip_if);
`endif // !`ifdef USE_VIP_SNPS
`ifdef USE_VIP_SNPS_APB
           uvm_config_db#(svt_apb_vif)::set(uvm_root::get(), 
            "", "vif", apb_vip_if);
`endif
    uvm_config_db#(virtual <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_apb_if)::set(.cntxt( uvm_root::get()),
                                        .inst_name( "" ),
                                        .field_name( "m_apb_if" ),
                                        .value(m_apb_if ));

   uvm_config_db#(virtual <%=obj.DiiInfo[obj.Id].strRtlNamePrefix%>_dii_rtl_if)::set(.cntxt( null ),
                                        .inst_name( "uvm_test_top" ),
                                        .field_name( "m_dii_rtl_if" ),
                                        .value( m_dii_rtl_if ));

    uvm_config_db#(virtual <%=obj.BlockId%>_q_chnl_if )::set(.cntxt( uvm_root::get()),
                                        .inst_name( "" ),
                                        .field_name( "m_q_chnl_if" ),
                                        .value(m_q_chnl_if ));



    system_quiesce = new("system_quiesce");
    system_unquiesce = new("system_unquiesce");


    uvm_config_db#(uvm_event)::set(.cntxt(null),
                                        .inst_name( "uvm_test_top.m_env" ),
                                        .field_name( "system_quiesce" ),
                                        .value( system_quiesce));
    uvm_config_db#(uvm_event)::set(.cntxt(null),
                                        .inst_name( "uvm_test_top.m_env" ),
                                        .field_name( "system_unquiesce" ),
                                        .value( system_unquiesce));



    injectSingleErrRtt = new("injectSingleErrRtt");
    injectDoubleErrRtt = new("injectDoubleErrRtt");


    checkCELR = new("checkCELR");
    checkUELR = new("checkUELR");


    forceClkgate   = new("forceClkgate");
    releaseClkgate = new("releaseClkgate");


    uvm_config_db#(uvm_event)::set(.cntxt(null),
                                        .inst_name( "uvm_test_top.m_env" ),
                                        .field_name( "injectSingleErrRtt" ),
                                        .value( injectSingleErrRtt));
    uvm_config_db#(uvm_event)::set(.cntxt(null),
                                        .inst_name( "uvm_test_top.m_env" ),
                                        .field_name( "injectDoubleErrRtt" ),
                                        .value( injectDoubleErrRtt));

    uvm_config_db#(uvm_event)::set(.cntxt(null),
                                        .inst_name( "uvm_test_top.m_env" ),
                                        .field_name( "checkCELR" ),
                                        .value( checkCELR));
    uvm_config_db#(uvm_event)::set(.cntxt(null),
                                        .inst_name( "uvm_test_top.m_env" ),
                                        .field_name( "checkUELR" ),
                                        .value( checkUELR));

    uvm_config_db#(uvm_event)::set(.cntxt( uvm_root::get()),
                                        .inst_name( "" ),
                                        .field_name( "forceClkgate" ),
                                        .value(forceClkgate));

    uvm_config_db#(uvm_event)::set(.cntxt( uvm_root::get()),
                                        .inst_name( "" ),
                                        .field_name( "releaseClkgate" ),
                                        .value(releaseClkgate));


//`ifdef VCS_SIM,CDNS
`ifdef DUMP_ON
  if ($test$plusargs("en_dump")) begin
  `ifdef VCS
   $vcdpluson;
  `elsif CDNS
   $shm_open ( "waves.shm" ) ;
   $shm_probe ( "ACMS" ) ;
  `endif
  end
`endif


    //force m_smis to 0 which are not yet connected
    force m_smi0_rx_smi_if.smi_msg_err = 0;
    force m_smi1_rx_smi_if.smi_msg_err = 0;
    force m_smi2_rx_smi_if.smi_msg_err = 0;

 <% for (var i=0; i<obj.DiiInfo[obj.Id].interfaces.smiTxInt.length; i++) {%>
    //setup for rx interface ready not ready ranges
    m_smi<%=i%>_rx_smi_if.my_smi_rx_id = <%=i%>;
 <%}%>

  run_test("dii_test");
  $finish;

end

       assign u_csr_probe_if.IRQ_C     = tb_top.dut.<%=obj.DiiInfo[obj.Id].interfaces.irqInt.name%>c;
       assign u_csr_probe_if.IRQ_UC    = tb_top.dut.<%=obj.DiiInfo[obj.Id].interfaces.irqInt.name%>uc;
<% if(obj.useResiliency) { %>
       assign u_csr_probe_if.fault_mission_fault = tb_top.dut.fault_mission_fault;
       assign u_csr_probe_if.fault_latent_fault = tb_top.dut.fault_latent_fault;
       assign u_csr_probe_if.cerr_threshold          = tb_top.dut.u_dii_fault_checker.cerr_threshold;
       assign u_csr_probe_if.cerr_counter            = tb_top.dut.u_dii_fault_checker.cerr_counter;
       assign u_csr_probe_if.cerr_over_thres_fault   = tb_top.dut.u_dii_fault_checker.cerr_over_thres_fault;

<% } %>
        // sys_event timeout signals :

        assign u_csr_probe_if.timeout_threshold       = tb_top.dut.u_dii_unit.dii_csr.dii_csr_gen.DIIUTOCR_TimeOutThreshold_out;
        assign u_csr_probe_if.sys_timeout_threshold   = tb_top.dut.u_dii_unit.dii_csr.dii_csr_gen.DIIUSEPTOCR_TimeOutThreshold_out;
        assign u_csr_probe_if.uedr_timeout_err_det_en = tb_top.dut.u_dii_unit.dii_csr.dii_csr_gen.DIIUUEDR_TimeoutErrDetEn_out;
        assign u_csr_probe_if.uesr_errvld             = tb_top.dut.u_dii_unit.dii_csr.dii_csr_gen.DIIUUESR_ErrVld_out;
        assign u_csr_probe_if.uesr_err_type           = tb_top.dut.u_dii_unit.dii_csr.dii_csr_gen.DIIUUESR_ErrType_out;
        assign u_csr_probe_if.uesr_err_info           = tb_top.dut.u_dii_unit.dii_csr.dii_csr_gen.DIIUUESR_ErrInfo_out;
        //assign u_csr_probe_if.ueir_timeout_irq_en     = tb_top.dut.u_dii_unit.dii_csr.dii_csr_gen.DIIUUEIR_TimeoutErrIntEn_out;

        // Sys event signals :

        assign m_dii_rtl_if.event_in_req 		= tb_top.dut.u_dii_unit.u_sys_evt_coh_concerto.event_in_req;
        assign m_dii_rtl_if.event_in_ack 		= tb_top.dut.u_dii_unit.u_sys_evt_coh_concerto.event_in_ack;
        assign m_dii_rtl_if.event_err_valid 	= tb_top.dut.u_dii_unit.u_sys_evt_coh_concerto.csr_sys_evt_sender_err_vld;

        ////////////////
<% if(!obj.CUSTOMER_ENV) { %>
//Task calls end of simulation tasks and pending transaction methods
task assert_error(input string verbose, input string msg);
    uvm_component  m_comp[$];
    dii_scoreboard m_scb;

    $display(msg);
    $stacktrace;

    #1ns;  // give a chance for waveform dumping

    uvm_top.find_all("uvm_test_top.m_env.m_scb", m_comp, uvm_top);
    if(m_comp.size() == 0) begin
        `uvm_fatal("tb_top", "none of the components are found with specified name")
    end
    if(m_comp.size() > 1) begin
        foreach(m_comp[i]) 
            `uvm_info("tb_top", $psprintf("component: %s", m_comp[i].get_full_name()), UVM_LOW)
        `uvm_fatal("tb_top", "multiple components with same name are found, components are specified above")
    end

    if(verbose == "FATAL") begin 
        `uvm_fatal("assert_error", msg) 
    end else begin 
        `uvm_error("assert_error", msg) 
    end
endtask: assert_error
<% } %>


//Checking clock idle when qREQn and qACCEPTn are low (entered into pma)
<% if(obj.DiiInfo[obj.Id].usePma) { %>
assert_clk_idle_when_pma_asserted : assert property (
    @(posedge fr_clk) disable iff (!soft_rstn)
    (!m_q_chnl_if.QREQn && !m_q_chnl_if.QACCEPTn ) |-> !dut_clk
    ) else assert_error("ERROR", "Dut clock is not stable low when RTL entered into PMA");
<% } %>


endmodule
